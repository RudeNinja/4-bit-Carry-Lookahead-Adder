magic
tech scmos
timestamp 1638809964
<< nwell >>
rect -341 292 -243 324
rect -183 283 -54 302
rect -341 184 -287 216
rect -341 114 -243 146
rect -154 143 -92 166
rect -56 140 27 167
rect 56 117 185 136
rect -341 6 -287 38
rect -179 1 -117 24
rect -96 -13 -34 10
rect -341 -64 -243 -32
rect 3 -47 86 -20
rect 116 -44 245 -25
rect -188 -97 -126 -74
rect -98 -120 -15 -93
rect -341 -172 -287 -140
rect -341 -242 -243 -210
rect -160 -216 -98 -193
rect -77 -230 -15 -207
rect 6 -238 68 -215
rect 83 -283 166 -256
rect -341 -350 -287 -318
rect -145 -332 -83 -309
rect -62 -346 0 -323
rect 47 -400 130 -373
rect -147 -426 -85 -403
rect -54 -443 29 -416
<< ntransistor >>
rect -329 275 -327 285
rect -257 275 -255 285
rect -169 250 -167 259
rect -305 240 -303 250
rect -295 240 -293 250
rect -285 240 -283 250
rect -275 240 -273 250
rect -77 251 -75 260
rect -144 213 -142 223
rect -132 213 -130 223
rect -118 213 -116 223
rect -105 213 -103 223
rect -329 160 -327 170
rect -319 160 -317 170
rect -301 160 -299 170
rect -329 97 -327 107
rect -257 97 -255 107
rect -141 100 -139 108
rect -128 100 -126 108
rect -106 101 -104 109
rect -38 87 -36 95
rect -20 87 -18 95
rect 7 87 9 95
rect 70 84 72 93
rect -305 62 -303 72
rect -295 62 -293 72
rect -285 62 -283 72
rect -275 62 -273 72
rect 162 85 164 94
rect 95 47 97 57
rect 107 47 109 57
rect 121 47 123 57
rect 134 47 136 57
rect -329 -18 -327 -8
rect -319 -18 -317 -8
rect -301 -18 -299 -8
rect -166 -42 -164 -34
rect -153 -42 -151 -34
rect -131 -41 -129 -33
rect -83 -56 -81 -48
rect -70 -56 -68 -48
rect -48 -55 -46 -47
rect -329 -81 -327 -71
rect -257 -81 -255 -71
rect -305 -116 -303 -106
rect -295 -116 -293 -106
rect -285 -116 -283 -106
rect -275 -116 -273 -106
rect 130 -77 132 -68
rect 21 -100 23 -92
rect 39 -100 41 -92
rect 66 -100 68 -92
rect 222 -76 224 -67
rect -175 -140 -173 -132
rect -162 -140 -160 -132
rect -140 -139 -138 -131
rect 155 -114 157 -104
rect 167 -114 169 -104
rect 181 -114 183 -104
rect 194 -114 196 -104
rect -80 -173 -78 -165
rect -62 -173 -60 -165
rect -35 -173 -33 -165
rect -329 -196 -327 -186
rect -319 -196 -317 -186
rect -301 -196 -299 -186
rect -329 -259 -327 -249
rect -257 -259 -255 -249
rect -147 -259 -145 -251
rect -134 -259 -132 -251
rect -112 -258 -110 -250
rect -64 -273 -62 -265
rect -51 -273 -49 -265
rect -29 -272 -27 -264
rect 19 -281 21 -273
rect 32 -281 34 -273
rect 54 -280 56 -272
rect -305 -294 -303 -284
rect -295 -294 -293 -284
rect -285 -294 -283 -284
rect -275 -294 -273 -284
rect -329 -374 -327 -364
rect -319 -374 -317 -364
rect -301 -374 -299 -364
rect 101 -336 103 -328
rect 119 -336 121 -328
rect 146 -336 148 -328
rect -132 -375 -130 -367
rect -119 -375 -117 -367
rect -97 -374 -95 -366
rect -49 -389 -47 -381
rect -36 -389 -34 -381
rect -14 -388 -12 -380
rect -134 -469 -132 -461
rect -121 -469 -119 -461
rect -99 -468 -97 -460
rect 65 -453 67 -445
rect 83 -453 85 -445
rect 110 -453 112 -445
rect -36 -496 -34 -488
rect -18 -496 -16 -488
rect 9 -496 11 -488
<< ptransistor >>
rect -329 298 -327 318
rect -305 298 -303 318
rect -295 298 -293 318
rect -285 298 -283 318
rect -275 298 -273 318
rect -257 298 -255 318
rect -169 289 -167 296
rect -144 289 -142 296
rect -132 289 -130 296
rect -118 289 -116 296
rect -105 289 -103 296
rect -77 289 -75 296
rect -329 190 -327 210
rect -319 190 -317 210
rect -301 190 -299 210
rect -141 149 -139 160
rect -128 149 -126 160
rect -106 149 -104 160
rect -329 120 -327 140
rect -305 120 -303 140
rect -295 120 -293 140
rect -285 120 -283 140
rect -275 120 -273 140
rect -257 120 -255 140
rect -38 148 -36 159
rect -20 148 -18 159
rect 7 148 9 159
rect 70 123 72 130
rect 95 123 97 130
rect 107 123 109 130
rect 121 123 123 130
rect 134 123 136 130
rect 162 123 164 130
rect -329 12 -327 32
rect -319 12 -317 32
rect -301 12 -299 32
rect -166 7 -164 18
rect -153 7 -151 18
rect -131 7 -129 18
rect -83 -7 -81 4
rect -70 -7 -68 4
rect -48 -7 -46 4
rect -329 -58 -327 -38
rect -305 -58 -303 -38
rect -295 -58 -293 -38
rect -285 -58 -283 -38
rect -275 -58 -273 -38
rect -257 -58 -255 -38
rect 21 -39 23 -28
rect 39 -39 41 -28
rect 66 -39 68 -28
rect 130 -38 132 -31
rect 155 -38 157 -31
rect 167 -38 169 -31
rect 181 -38 183 -31
rect 194 -38 196 -31
rect 222 -38 224 -31
rect -175 -91 -173 -80
rect -162 -91 -160 -80
rect -140 -91 -138 -80
rect -80 -112 -78 -101
rect -62 -112 -60 -101
rect -35 -112 -33 -101
rect -329 -166 -327 -146
rect -319 -166 -317 -146
rect -301 -166 -299 -146
rect -147 -210 -145 -199
rect -134 -210 -132 -199
rect -112 -210 -110 -199
rect -329 -236 -327 -216
rect -305 -236 -303 -216
rect -295 -236 -293 -216
rect -285 -236 -283 -216
rect -275 -236 -273 -216
rect -257 -236 -255 -216
rect -64 -224 -62 -213
rect -51 -224 -49 -213
rect -29 -224 -27 -213
rect 19 -232 21 -221
rect 32 -232 34 -221
rect 54 -232 56 -221
rect 101 -275 103 -264
rect 119 -275 121 -264
rect 146 -275 148 -264
rect -329 -344 -327 -324
rect -319 -344 -317 -324
rect -301 -344 -299 -324
rect -132 -326 -130 -315
rect -119 -326 -117 -315
rect -97 -326 -95 -315
rect -49 -340 -47 -329
rect -36 -340 -34 -329
rect -14 -340 -12 -329
rect 65 -392 67 -381
rect 83 -392 85 -381
rect 110 -392 112 -381
rect -134 -420 -132 -409
rect -121 -420 -119 -409
rect -99 -420 -97 -409
rect -36 -435 -34 -424
rect -18 -435 -16 -424
rect 9 -435 11 -424
<< ndiffusion >>
rect -331 275 -329 285
rect -327 275 -325 285
rect -259 275 -257 285
rect -255 275 -253 285
rect -172 250 -169 259
rect -167 250 -164 259
rect -307 240 -305 250
rect -303 240 -301 250
rect -297 240 -295 250
rect -293 240 -291 250
rect -287 240 -285 250
rect -283 240 -281 250
rect -277 240 -275 250
rect -273 240 -271 250
rect -80 251 -77 260
rect -75 251 -72 260
rect -147 213 -144 223
rect -142 213 -139 223
rect -135 213 -132 223
rect -130 213 -127 223
rect -122 213 -118 223
rect -116 213 -113 223
rect -109 213 -105 223
rect -103 213 -100 223
rect -95 213 -93 223
rect -331 160 -329 170
rect -327 160 -319 170
rect -317 160 -315 170
rect -303 160 -301 170
rect -299 160 -297 170
rect -331 97 -329 107
rect -327 97 -325 107
rect -259 97 -257 107
rect -255 97 -253 107
rect -143 100 -141 108
rect -139 100 -128 108
rect -126 100 -125 108
rect -107 101 -106 109
rect -104 101 -102 109
rect -40 87 -38 95
rect -36 87 -30 95
rect -25 87 -20 95
rect -18 87 -14 95
rect 6 87 7 95
rect 9 87 12 95
rect 67 84 70 93
rect 72 84 75 93
rect -307 62 -305 72
rect -303 62 -301 72
rect -297 62 -295 72
rect -293 62 -291 72
rect -287 62 -285 72
rect -283 62 -281 72
rect -277 62 -275 72
rect -273 62 -271 72
rect 159 85 162 94
rect 164 85 167 94
rect 92 47 95 57
rect 97 47 100 57
rect 104 47 107 57
rect 109 47 112 57
rect 117 47 121 57
rect 123 47 126 57
rect 130 47 134 57
rect 136 47 139 57
rect 144 47 146 57
rect -331 -18 -329 -8
rect -327 -18 -319 -8
rect -317 -18 -315 -8
rect -303 -18 -301 -8
rect -299 -18 -297 -8
rect -168 -42 -166 -34
rect -164 -42 -153 -34
rect -151 -42 -150 -34
rect -132 -41 -131 -33
rect -129 -41 -127 -33
rect -85 -56 -83 -48
rect -81 -56 -70 -48
rect -68 -56 -67 -48
rect -49 -55 -48 -47
rect -46 -55 -44 -47
rect -331 -81 -329 -71
rect -327 -81 -325 -71
rect -259 -81 -257 -71
rect -255 -81 -253 -71
rect -307 -116 -305 -106
rect -303 -116 -301 -106
rect -297 -116 -295 -106
rect -293 -116 -291 -106
rect -287 -116 -285 -106
rect -283 -116 -281 -106
rect -277 -116 -275 -106
rect -273 -116 -271 -106
rect 127 -77 130 -68
rect 132 -77 135 -68
rect 19 -100 21 -92
rect 23 -100 29 -92
rect 34 -100 39 -92
rect 41 -100 45 -92
rect 65 -100 66 -92
rect 68 -100 71 -92
rect 219 -76 222 -67
rect 224 -76 227 -67
rect -177 -140 -175 -132
rect -173 -140 -162 -132
rect -160 -140 -159 -132
rect -141 -139 -140 -131
rect -138 -139 -136 -131
rect 152 -114 155 -104
rect 157 -114 160 -104
rect 164 -114 167 -104
rect 169 -114 172 -104
rect 177 -114 181 -104
rect 183 -114 186 -104
rect 190 -114 194 -104
rect 196 -114 199 -104
rect 204 -114 206 -104
rect -82 -173 -80 -165
rect -78 -173 -72 -165
rect -67 -173 -62 -165
rect -60 -173 -56 -165
rect -36 -173 -35 -165
rect -33 -173 -30 -165
rect -331 -196 -329 -186
rect -327 -196 -319 -186
rect -317 -196 -315 -186
rect -303 -196 -301 -186
rect -299 -196 -297 -186
rect -331 -259 -329 -249
rect -327 -259 -325 -249
rect -259 -259 -257 -249
rect -255 -259 -253 -249
rect -149 -259 -147 -251
rect -145 -259 -134 -251
rect -132 -259 -131 -251
rect -113 -258 -112 -250
rect -110 -258 -108 -250
rect -66 -273 -64 -265
rect -62 -273 -51 -265
rect -49 -273 -48 -265
rect -30 -272 -29 -264
rect -27 -272 -25 -264
rect 17 -281 19 -273
rect 21 -281 32 -273
rect 34 -281 35 -273
rect 53 -280 54 -272
rect 56 -280 58 -272
rect -307 -294 -305 -284
rect -303 -294 -301 -284
rect -297 -294 -295 -284
rect -293 -294 -291 -284
rect -287 -294 -285 -284
rect -283 -294 -281 -284
rect -277 -294 -275 -284
rect -273 -294 -271 -284
rect -331 -374 -329 -364
rect -327 -374 -319 -364
rect -317 -374 -315 -364
rect -303 -374 -301 -364
rect -299 -374 -297 -364
rect 99 -336 101 -328
rect 103 -336 109 -328
rect 114 -336 119 -328
rect 121 -336 125 -328
rect 145 -336 146 -328
rect 148 -336 151 -328
rect -134 -375 -132 -367
rect -130 -375 -119 -367
rect -117 -375 -116 -367
rect -98 -374 -97 -366
rect -95 -374 -93 -366
rect -51 -389 -49 -381
rect -47 -389 -36 -381
rect -34 -389 -33 -381
rect -15 -388 -14 -380
rect -12 -388 -10 -380
rect -136 -469 -134 -461
rect -132 -469 -121 -461
rect -119 -469 -118 -461
rect -100 -468 -99 -460
rect -97 -468 -95 -460
rect 63 -453 65 -445
rect 67 -453 73 -445
rect 78 -453 83 -445
rect 85 -453 89 -445
rect 109 -453 110 -445
rect 112 -453 115 -445
rect -38 -496 -36 -488
rect -34 -496 -28 -488
rect -23 -496 -18 -488
rect -16 -496 -12 -488
rect 8 -496 9 -488
rect 11 -496 14 -488
<< pdiffusion >>
rect -331 298 -329 318
rect -327 298 -325 318
rect -307 298 -305 318
rect -303 298 -295 318
rect -293 298 -291 318
rect -287 298 -285 318
rect -283 298 -275 318
rect -273 298 -271 318
rect -259 298 -257 318
rect -255 298 -253 318
rect -172 289 -169 296
rect -167 289 -164 296
rect -147 289 -144 296
rect -142 289 -132 296
rect -130 289 -126 296
rect -122 289 -118 296
rect -116 289 -105 296
rect -103 289 -98 296
rect -80 289 -77 296
rect -75 289 -72 296
rect -331 190 -329 210
rect -327 190 -325 210
rect -321 190 -319 210
rect -317 190 -315 210
rect -303 190 -301 210
rect -299 190 -297 210
rect -143 149 -141 160
rect -139 149 -133 160
rect -129 149 -128 160
rect -126 149 -124 160
rect -110 149 -106 160
rect -104 149 -102 160
rect -331 120 -329 140
rect -327 120 -325 140
rect -307 120 -305 140
rect -303 120 -295 140
rect -293 120 -291 140
rect -287 120 -285 140
rect -283 120 -275 140
rect -273 120 -271 140
rect -259 120 -257 140
rect -255 120 -253 140
rect -42 148 -38 159
rect -36 148 -20 159
rect -18 148 -14 159
rect -4 148 -1 159
rect 4 148 7 159
rect 9 148 12 159
rect 16 148 18 159
rect 67 123 70 130
rect 72 123 75 130
rect 92 123 95 130
rect 97 123 107 130
rect 109 123 113 130
rect 117 123 121 130
rect 123 123 134 130
rect 136 123 141 130
rect 159 123 162 130
rect 164 123 167 130
rect -331 12 -329 32
rect -327 12 -325 32
rect -321 12 -319 32
rect -317 12 -315 32
rect -303 12 -301 32
rect -299 12 -297 32
rect -168 7 -166 18
rect -164 7 -158 18
rect -154 7 -153 18
rect -151 7 -149 18
rect -135 7 -131 18
rect -129 7 -127 18
rect -85 -7 -83 4
rect -81 -7 -75 4
rect -71 -7 -70 4
rect -68 -7 -66 4
rect -52 -7 -48 4
rect -46 -7 -44 4
rect -331 -58 -329 -38
rect -327 -58 -325 -38
rect -307 -58 -305 -38
rect -303 -58 -295 -38
rect -293 -58 -291 -38
rect -287 -58 -285 -38
rect -283 -58 -275 -38
rect -273 -58 -271 -38
rect -259 -58 -257 -38
rect -255 -58 -253 -38
rect 17 -39 21 -28
rect 23 -39 39 -28
rect 41 -39 45 -28
rect 55 -39 58 -28
rect 63 -39 66 -28
rect 68 -39 71 -28
rect 75 -39 77 -28
rect 127 -38 130 -31
rect 132 -38 135 -31
rect 152 -38 155 -31
rect 157 -38 167 -31
rect 169 -38 173 -31
rect 177 -38 181 -31
rect 183 -38 194 -31
rect 196 -38 201 -31
rect 219 -38 222 -31
rect 224 -38 227 -31
rect -177 -91 -175 -80
rect -173 -91 -167 -80
rect -163 -91 -162 -80
rect -160 -91 -158 -80
rect -144 -91 -140 -80
rect -138 -91 -136 -80
rect -84 -112 -80 -101
rect -78 -112 -62 -101
rect -60 -112 -56 -101
rect -46 -112 -43 -101
rect -38 -112 -35 -101
rect -33 -112 -30 -101
rect -26 -112 -24 -101
rect -331 -166 -329 -146
rect -327 -166 -325 -146
rect -321 -166 -319 -146
rect -317 -166 -315 -146
rect -303 -166 -301 -146
rect -299 -166 -297 -146
rect -149 -210 -147 -199
rect -145 -210 -139 -199
rect -135 -210 -134 -199
rect -132 -210 -130 -199
rect -116 -210 -112 -199
rect -110 -210 -108 -199
rect -331 -236 -329 -216
rect -327 -236 -325 -216
rect -307 -236 -305 -216
rect -303 -236 -295 -216
rect -293 -236 -291 -216
rect -287 -236 -285 -216
rect -283 -236 -275 -216
rect -273 -236 -271 -216
rect -259 -236 -257 -216
rect -255 -236 -253 -216
rect -66 -224 -64 -213
rect -62 -224 -56 -213
rect -52 -224 -51 -213
rect -49 -224 -47 -213
rect -33 -224 -29 -213
rect -27 -224 -25 -213
rect 17 -232 19 -221
rect 21 -232 27 -221
rect 31 -232 32 -221
rect 34 -232 36 -221
rect 50 -232 54 -221
rect 56 -232 58 -221
rect 97 -275 101 -264
rect 103 -275 119 -264
rect 121 -275 125 -264
rect 135 -275 138 -264
rect 143 -275 146 -264
rect 148 -275 151 -264
rect 155 -275 157 -264
rect -331 -344 -329 -324
rect -327 -344 -325 -324
rect -321 -344 -319 -324
rect -317 -344 -315 -324
rect -303 -344 -301 -324
rect -299 -344 -297 -324
rect -134 -326 -132 -315
rect -130 -326 -124 -315
rect -120 -326 -119 -315
rect -117 -326 -115 -315
rect -101 -326 -97 -315
rect -95 -326 -93 -315
rect -51 -340 -49 -329
rect -47 -340 -41 -329
rect -37 -340 -36 -329
rect -34 -340 -32 -329
rect -18 -340 -14 -329
rect -12 -340 -10 -329
rect 61 -392 65 -381
rect 67 -392 83 -381
rect 85 -392 89 -381
rect 99 -392 102 -381
rect 107 -392 110 -381
rect 112 -392 115 -381
rect 119 -392 121 -381
rect -136 -420 -134 -409
rect -132 -420 -126 -409
rect -122 -420 -121 -409
rect -119 -420 -117 -409
rect -103 -420 -99 -409
rect -97 -420 -95 -409
rect -40 -435 -36 -424
rect -34 -435 -18 -424
rect -16 -435 -12 -424
rect -2 -435 1 -424
rect 6 -435 9 -424
rect 11 -435 14 -424
rect 18 -435 20 -424
<< ndcontact >>
rect -335 275 -331 285
rect -325 275 -321 285
rect -263 275 -259 285
rect -253 275 -249 285
rect -176 250 -172 259
rect -164 250 -160 259
rect -311 240 -307 250
rect -301 240 -297 250
rect -291 240 -287 250
rect -281 240 -277 250
rect -271 240 -267 250
rect -84 251 -80 260
rect -72 251 -68 260
rect -152 213 -147 223
rect -139 213 -135 223
rect -127 213 -122 223
rect -113 213 -109 223
rect -100 213 -95 223
rect -335 160 -331 170
rect -315 160 -311 170
rect -307 160 -303 170
rect -297 160 -293 170
rect -335 97 -331 107
rect -325 97 -321 107
rect -263 97 -259 107
rect -253 97 -249 107
rect -147 100 -143 108
rect -125 100 -121 108
rect -111 101 -107 109
rect -102 101 -98 109
rect -45 87 -40 95
rect -30 87 -25 95
rect -14 87 -9 95
rect 1 87 6 95
rect 12 87 16 95
rect 63 84 67 93
rect 75 84 79 93
rect -311 62 -307 72
rect -301 62 -297 72
rect -291 62 -287 72
rect -281 62 -277 72
rect -271 62 -267 72
rect 155 85 159 94
rect 167 85 171 94
rect 87 47 92 57
rect 100 47 104 57
rect 112 47 117 57
rect 126 47 130 57
rect 139 47 144 57
rect -335 -18 -331 -8
rect -315 -18 -311 -8
rect -307 -18 -303 -8
rect -297 -18 -293 -8
rect -172 -42 -168 -34
rect -150 -42 -146 -34
rect -136 -41 -132 -33
rect -127 -41 -123 -33
rect -89 -56 -85 -48
rect -67 -56 -63 -48
rect -53 -55 -49 -47
rect -44 -55 -40 -47
rect -335 -81 -331 -71
rect -325 -81 -321 -71
rect -263 -81 -259 -71
rect -253 -81 -249 -71
rect -311 -116 -307 -106
rect -301 -116 -297 -106
rect -291 -116 -287 -106
rect -281 -116 -277 -106
rect -271 -116 -267 -106
rect 123 -77 127 -68
rect 135 -77 139 -68
rect 14 -100 19 -92
rect 29 -100 34 -92
rect 45 -100 50 -92
rect 60 -100 65 -92
rect 71 -100 75 -92
rect 215 -76 219 -67
rect 227 -76 231 -67
rect -181 -140 -177 -132
rect -159 -140 -155 -132
rect -145 -139 -141 -131
rect -136 -139 -132 -131
rect 147 -114 152 -104
rect 160 -114 164 -104
rect 172 -114 177 -104
rect 186 -114 190 -104
rect 199 -114 204 -104
rect -87 -173 -82 -165
rect -72 -173 -67 -165
rect -56 -173 -51 -165
rect -41 -173 -36 -165
rect -30 -173 -26 -165
rect -335 -196 -331 -186
rect -315 -196 -311 -186
rect -307 -196 -303 -186
rect -297 -196 -293 -186
rect -335 -259 -331 -249
rect -325 -259 -321 -249
rect -263 -259 -259 -249
rect -253 -259 -249 -249
rect -153 -259 -149 -251
rect -131 -259 -127 -251
rect -117 -258 -113 -250
rect -108 -258 -104 -250
rect -70 -273 -66 -265
rect -48 -273 -44 -265
rect -34 -272 -30 -264
rect -25 -272 -21 -264
rect 13 -281 17 -273
rect 35 -281 39 -273
rect 49 -280 53 -272
rect 58 -280 62 -272
rect -311 -294 -307 -284
rect -301 -294 -297 -284
rect -291 -294 -287 -284
rect -281 -294 -277 -284
rect -271 -294 -267 -284
rect -335 -374 -331 -364
rect -315 -374 -311 -364
rect -307 -374 -303 -364
rect -297 -374 -293 -364
rect 94 -336 99 -328
rect 109 -336 114 -328
rect 125 -336 130 -328
rect 140 -336 145 -328
rect 151 -336 155 -328
rect -138 -375 -134 -367
rect -116 -375 -112 -367
rect -102 -374 -98 -366
rect -93 -374 -89 -366
rect -55 -389 -51 -381
rect -33 -389 -29 -381
rect -19 -388 -15 -380
rect -10 -388 -6 -380
rect -140 -469 -136 -461
rect -118 -469 -114 -461
rect -104 -468 -100 -460
rect -95 -468 -91 -460
rect 58 -453 63 -445
rect 73 -453 78 -445
rect 89 -453 94 -445
rect 104 -453 109 -445
rect 115 -453 119 -445
rect -43 -496 -38 -488
rect -28 -496 -23 -488
rect -12 -496 -7 -488
rect 3 -496 8 -488
rect 14 -496 18 -488
<< pdcontact >>
rect -335 298 -331 318
rect -325 298 -321 318
rect -311 298 -307 318
rect -291 298 -287 318
rect -271 298 -267 318
rect -263 298 -259 318
rect -253 298 -249 318
rect -176 289 -172 296
rect -164 289 -160 296
rect -151 289 -147 296
rect -126 289 -122 296
rect -98 289 -94 296
rect -84 289 -80 296
rect -72 289 -68 296
rect -335 190 -331 210
rect -325 190 -321 210
rect -315 190 -311 210
rect -307 190 -303 210
rect -297 190 -293 210
rect -148 149 -143 160
rect -133 149 -129 160
rect -124 149 -120 160
rect -114 149 -110 160
rect -102 149 -98 160
rect -335 120 -331 140
rect -325 120 -321 140
rect -311 120 -307 140
rect -291 120 -287 140
rect -271 120 -267 140
rect -263 120 -259 140
rect -253 120 -249 140
rect -48 148 -42 159
rect -14 148 -9 159
rect -1 148 4 159
rect 12 148 16 159
rect 63 123 67 130
rect 75 123 79 130
rect 88 123 92 130
rect 113 123 117 130
rect 141 123 145 130
rect 155 123 159 130
rect 167 123 171 130
rect -335 12 -331 32
rect -325 12 -321 32
rect -315 12 -311 32
rect -307 12 -303 32
rect -297 12 -293 32
rect -173 7 -168 18
rect -158 7 -154 18
rect -149 7 -145 18
rect -139 7 -135 18
rect -127 7 -123 18
rect -90 -7 -85 4
rect -75 -7 -71 4
rect -66 -7 -62 4
rect -56 -7 -52 4
rect -44 -7 -40 4
rect -335 -58 -331 -38
rect -325 -58 -321 -38
rect -311 -58 -307 -38
rect -291 -58 -287 -38
rect -271 -58 -267 -38
rect -263 -58 -259 -38
rect -253 -58 -249 -38
rect 11 -39 17 -28
rect 45 -39 50 -28
rect 58 -39 63 -28
rect 71 -39 75 -28
rect 123 -38 127 -31
rect 135 -38 139 -31
rect 148 -38 152 -31
rect 173 -38 177 -31
rect 201 -38 205 -31
rect 215 -38 219 -31
rect 227 -38 231 -31
rect -182 -91 -177 -80
rect -167 -91 -163 -80
rect -158 -91 -154 -80
rect -148 -91 -144 -80
rect -136 -91 -132 -80
rect -90 -112 -84 -101
rect -56 -112 -51 -101
rect -43 -112 -38 -101
rect -30 -112 -26 -101
rect -335 -166 -331 -146
rect -325 -166 -321 -146
rect -315 -166 -311 -146
rect -307 -166 -303 -146
rect -297 -166 -293 -146
rect -154 -210 -149 -199
rect -139 -210 -135 -199
rect -130 -210 -126 -199
rect -120 -210 -116 -199
rect -108 -210 -104 -199
rect -335 -236 -331 -216
rect -325 -236 -321 -216
rect -311 -236 -307 -216
rect -291 -236 -287 -216
rect -271 -236 -267 -216
rect -263 -236 -259 -216
rect -253 -236 -249 -216
rect -71 -224 -66 -213
rect -56 -224 -52 -213
rect -47 -224 -43 -213
rect -37 -224 -33 -213
rect -25 -224 -21 -213
rect 12 -232 17 -221
rect 27 -232 31 -221
rect 36 -232 40 -221
rect 46 -232 50 -221
rect 58 -232 62 -221
rect 91 -275 97 -264
rect 125 -275 130 -264
rect 138 -275 143 -264
rect 151 -275 155 -264
rect -335 -344 -331 -324
rect -325 -344 -321 -324
rect -315 -344 -311 -324
rect -307 -344 -303 -324
rect -297 -344 -293 -324
rect -139 -326 -134 -315
rect -124 -326 -120 -315
rect -115 -326 -111 -315
rect -105 -326 -101 -315
rect -93 -326 -89 -315
rect -56 -340 -51 -329
rect -41 -340 -37 -329
rect -32 -340 -28 -329
rect -22 -340 -18 -329
rect -10 -340 -6 -329
rect 55 -392 61 -381
rect 89 -392 94 -381
rect 102 -392 107 -381
rect 115 -392 119 -381
rect -141 -420 -136 -409
rect -126 -420 -122 -409
rect -117 -420 -113 -409
rect -107 -420 -103 -409
rect -95 -420 -91 -409
rect -46 -435 -40 -424
rect -12 -435 -7 -424
rect 1 -435 6 -424
rect 14 -435 18 -424
<< polysilicon >>
rect -329 318 -327 321
rect -305 318 -303 321
rect -295 318 -293 321
rect -285 318 -283 321
rect -275 318 -273 321
rect -257 318 -255 321
rect -329 285 -327 298
rect -329 272 -327 275
rect -305 250 -303 298
rect -295 250 -293 298
rect -285 250 -283 298
rect -275 250 -273 298
rect -257 285 -255 298
rect -169 296 -167 299
rect -144 296 -142 299
rect -132 296 -130 299
rect -118 296 -116 299
rect -105 296 -103 299
rect -77 296 -75 299
rect -257 272 -255 275
rect -169 259 -167 289
rect -169 247 -167 250
rect -305 237 -303 240
rect -295 237 -293 240
rect -285 237 -283 240
rect -275 237 -273 240
rect -144 223 -142 289
rect -132 223 -130 289
rect -118 223 -116 289
rect -105 223 -103 289
rect -77 260 -75 289
rect -77 247 -75 251
rect -329 210 -327 213
rect -319 210 -317 213
rect -301 210 -299 213
rect -144 210 -142 213
rect -132 210 -130 213
rect -118 210 -116 213
rect -105 210 -103 213
rect -329 170 -327 190
rect -319 170 -317 190
rect -301 170 -299 190
rect -141 160 -139 163
rect -128 160 -126 163
rect -106 160 -104 163
rect -329 157 -327 160
rect -319 157 -317 160
rect -301 157 -299 160
rect -38 159 -36 163
rect -20 159 -18 163
rect 7 159 9 162
rect -329 140 -327 143
rect -305 140 -303 143
rect -295 140 -293 143
rect -285 140 -283 143
rect -275 140 -273 143
rect -257 140 -255 143
rect -329 107 -327 120
rect -329 94 -327 97
rect -305 72 -303 120
rect -295 72 -293 120
rect -285 72 -283 120
rect -275 72 -273 120
rect -257 107 -255 120
rect -141 108 -139 149
rect -128 108 -126 149
rect -106 109 -104 149
rect -141 97 -139 100
rect -128 97 -126 100
rect -106 98 -104 101
rect -257 94 -255 97
rect -38 95 -36 148
rect -20 95 -18 148
rect 7 95 9 148
rect 70 130 72 133
rect 95 130 97 133
rect 107 130 109 133
rect 121 130 123 133
rect 134 130 136 133
rect 162 130 164 133
rect 70 93 72 123
rect -38 84 -36 87
rect -20 84 -18 87
rect 7 84 9 87
rect 70 81 72 84
rect -305 59 -303 62
rect -295 59 -293 62
rect -285 59 -283 62
rect -275 59 -273 62
rect 95 57 97 123
rect 107 57 109 123
rect 121 57 123 123
rect 134 57 136 123
rect 162 94 164 123
rect 162 81 164 85
rect 95 44 97 47
rect 107 44 109 47
rect 121 44 123 47
rect 134 44 136 47
rect -329 32 -327 35
rect -319 32 -317 35
rect -301 32 -299 35
rect -166 18 -164 21
rect -153 18 -151 21
rect -131 18 -129 21
rect -329 -8 -327 12
rect -319 -8 -317 12
rect -301 -8 -299 12
rect -329 -21 -327 -18
rect -319 -21 -317 -18
rect -301 -21 -299 -18
rect -166 -34 -164 7
rect -153 -34 -151 7
rect -131 -33 -129 7
rect -83 4 -81 7
rect -70 4 -68 7
rect -48 4 -46 7
rect -329 -38 -327 -35
rect -305 -38 -303 -35
rect -295 -38 -293 -35
rect -285 -38 -283 -35
rect -275 -38 -273 -35
rect -257 -38 -255 -35
rect -166 -45 -164 -42
rect -153 -45 -151 -42
rect -131 -44 -129 -41
rect -83 -48 -81 -7
rect -70 -48 -68 -7
rect -48 -47 -46 -7
rect 21 -28 23 -24
rect 39 -28 41 -24
rect 66 -28 68 -25
rect 130 -31 132 -28
rect 155 -31 157 -28
rect 167 -31 169 -28
rect 181 -31 183 -28
rect 194 -31 196 -28
rect 222 -31 224 -28
rect -329 -71 -327 -58
rect -329 -84 -327 -81
rect -305 -106 -303 -58
rect -295 -106 -293 -58
rect -285 -106 -283 -58
rect -275 -106 -273 -58
rect -257 -71 -255 -58
rect -83 -59 -81 -56
rect -70 -59 -68 -56
rect -48 -58 -46 -55
rect -175 -80 -173 -77
rect -162 -80 -160 -77
rect -140 -80 -138 -77
rect -257 -84 -255 -81
rect -305 -119 -303 -116
rect -295 -119 -293 -116
rect -285 -119 -283 -116
rect -275 -119 -273 -116
rect -175 -132 -173 -91
rect -162 -132 -160 -91
rect -140 -131 -138 -91
rect 21 -92 23 -39
rect 39 -92 41 -39
rect 66 -92 68 -39
rect 130 -68 132 -38
rect 130 -80 132 -77
rect -80 -101 -78 -97
rect -62 -101 -60 -97
rect -35 -101 -33 -98
rect 21 -103 23 -100
rect 39 -103 41 -100
rect 66 -103 68 -100
rect 155 -104 157 -38
rect 167 -104 169 -38
rect 181 -104 183 -38
rect 194 -104 196 -38
rect 222 -67 224 -38
rect 222 -80 224 -76
rect -175 -143 -173 -140
rect -162 -143 -160 -140
rect -140 -142 -138 -139
rect -329 -146 -327 -143
rect -319 -146 -317 -143
rect -301 -146 -299 -143
rect -80 -165 -78 -112
rect -62 -165 -60 -112
rect -35 -165 -33 -112
rect 155 -117 157 -114
rect 167 -117 169 -114
rect 181 -117 183 -114
rect 194 -117 196 -114
rect -329 -186 -327 -166
rect -319 -186 -317 -166
rect -301 -186 -299 -166
rect -80 -176 -78 -173
rect -62 -176 -60 -173
rect -35 -176 -33 -173
rect -329 -199 -327 -196
rect -319 -199 -317 -196
rect -301 -199 -299 -196
rect -147 -199 -145 -196
rect -134 -199 -132 -196
rect -112 -199 -110 -196
rect -329 -216 -327 -213
rect -305 -216 -303 -213
rect -295 -216 -293 -213
rect -285 -216 -283 -213
rect -275 -216 -273 -213
rect -257 -216 -255 -213
rect -329 -249 -327 -236
rect -329 -262 -327 -259
rect -305 -284 -303 -236
rect -295 -284 -293 -236
rect -285 -284 -283 -236
rect -275 -284 -273 -236
rect -257 -249 -255 -236
rect -147 -251 -145 -210
rect -134 -251 -132 -210
rect -112 -250 -110 -210
rect -64 -213 -62 -210
rect -51 -213 -49 -210
rect -29 -213 -27 -210
rect 19 -221 21 -218
rect 32 -221 34 -218
rect 54 -221 56 -218
rect -257 -262 -255 -259
rect -147 -262 -145 -259
rect -134 -262 -132 -259
rect -112 -261 -110 -258
rect -64 -265 -62 -224
rect -51 -265 -49 -224
rect -29 -264 -27 -224
rect -64 -276 -62 -273
rect -51 -276 -49 -273
rect -29 -275 -27 -272
rect 19 -273 21 -232
rect 32 -273 34 -232
rect 54 -272 56 -232
rect 101 -264 103 -260
rect 119 -264 121 -260
rect 146 -264 148 -261
rect 19 -284 21 -281
rect 32 -284 34 -281
rect 54 -283 56 -280
rect -305 -297 -303 -294
rect -295 -297 -293 -294
rect -285 -297 -283 -294
rect -275 -297 -273 -294
rect -132 -315 -130 -312
rect -119 -315 -117 -312
rect -97 -315 -95 -312
rect -329 -324 -327 -321
rect -319 -324 -317 -321
rect -301 -324 -299 -321
rect -329 -364 -327 -344
rect -319 -364 -317 -344
rect -301 -364 -299 -344
rect -132 -367 -130 -326
rect -119 -367 -117 -326
rect -97 -366 -95 -326
rect -49 -329 -47 -326
rect -36 -329 -34 -326
rect -14 -329 -12 -326
rect 101 -328 103 -275
rect 119 -328 121 -275
rect 146 -328 148 -275
rect 101 -339 103 -336
rect 119 -339 121 -336
rect 146 -339 148 -336
rect -329 -377 -327 -374
rect -319 -377 -317 -374
rect -301 -377 -299 -374
rect -132 -378 -130 -375
rect -119 -378 -117 -375
rect -97 -377 -95 -374
rect -49 -381 -47 -340
rect -36 -381 -34 -340
rect -14 -380 -12 -340
rect 65 -381 67 -377
rect 83 -381 85 -377
rect 110 -381 112 -378
rect -49 -392 -47 -389
rect -36 -392 -34 -389
rect -14 -391 -12 -388
rect -134 -409 -132 -406
rect -121 -409 -119 -406
rect -99 -409 -97 -406
rect -134 -461 -132 -420
rect -121 -461 -119 -420
rect -99 -460 -97 -420
rect -36 -424 -34 -420
rect -18 -424 -16 -420
rect 9 -424 11 -421
rect -134 -472 -132 -469
rect -121 -472 -119 -469
rect -99 -471 -97 -468
rect -36 -488 -34 -435
rect -18 -488 -16 -435
rect 9 -488 11 -435
rect 65 -445 67 -392
rect 83 -445 85 -392
rect 110 -445 112 -392
rect 65 -456 67 -453
rect 83 -456 85 -453
rect 110 -456 112 -453
rect -36 -499 -34 -496
rect -18 -499 -16 -496
rect 9 -499 11 -496
<< polycontact >>
rect -333 288 -329 292
rect -309 256 -305 260
rect -299 288 -295 292
rect -289 267 -285 271
rect -273 285 -269 289
rect -255 288 -251 292
rect -173 269 -169 273
rect -148 229 -144 233
rect -136 267 -132 271
rect -122 255 -118 259
rect -103 267 -99 271
rect -75 267 -71 271
rect -333 180 -329 184
rect -323 173 -319 177
rect -305 173 -301 177
rect -145 134 -141 138
rect -333 110 -329 114
rect -309 78 -305 82
rect -299 110 -295 114
rect -289 89 -285 93
rect -273 107 -269 111
rect -255 110 -251 114
rect -132 117 -128 121
rect -110 132 -106 136
rect -43 132 -38 137
rect -25 118 -20 123
rect 3 129 7 134
rect 66 103 70 107
rect 91 63 95 67
rect 103 101 107 105
rect 117 89 121 93
rect 136 101 140 105
rect 164 101 168 105
rect -333 2 -329 6
rect -323 -5 -319 -1
rect -305 -5 -301 -1
rect -170 -8 -166 -4
rect -157 -25 -153 -21
rect -135 -10 -131 -6
rect -87 -22 -83 -18
rect -74 -39 -70 -35
rect -52 -24 -48 -20
rect 16 -55 21 -50
rect -333 -68 -329 -64
rect -309 -100 -305 -96
rect -299 -68 -295 -64
rect -289 -89 -285 -85
rect -273 -71 -269 -67
rect -255 -68 -251 -64
rect -179 -106 -175 -102
rect -166 -123 -162 -119
rect -144 -108 -140 -104
rect 34 -69 39 -64
rect 62 -58 66 -53
rect 126 -58 130 -54
rect 151 -98 155 -94
rect 163 -60 167 -56
rect 177 -72 181 -68
rect 196 -60 200 -56
rect 224 -60 228 -56
rect -85 -128 -80 -123
rect -67 -142 -62 -137
rect -39 -131 -35 -126
rect -333 -176 -329 -172
rect -323 -183 -319 -179
rect -305 -183 -301 -179
rect -151 -225 -147 -221
rect -333 -246 -329 -242
rect -309 -278 -305 -274
rect -299 -246 -295 -242
rect -289 -267 -285 -263
rect -273 -249 -269 -245
rect -255 -246 -251 -242
rect -138 -242 -134 -238
rect -116 -227 -112 -223
rect -68 -239 -64 -235
rect -55 -256 -51 -252
rect -33 -241 -29 -237
rect 15 -247 19 -243
rect 28 -264 32 -260
rect 50 -249 54 -245
rect 96 -291 101 -286
rect -136 -341 -132 -337
rect -333 -354 -329 -350
rect -323 -361 -319 -357
rect -305 -361 -301 -357
rect -123 -358 -119 -354
rect -101 -343 -97 -339
rect 114 -305 119 -300
rect 142 -294 146 -289
rect -53 -355 -49 -351
rect -40 -372 -36 -368
rect -18 -357 -14 -353
rect 60 -408 65 -403
rect -138 -435 -134 -431
rect -125 -452 -121 -448
rect -103 -437 -99 -433
rect -41 -451 -36 -446
rect -23 -465 -18 -460
rect 5 -454 9 -449
rect 78 -422 83 -417
rect 106 -411 110 -406
<< metal1 >>
rect -341 321 -243 325
rect -335 318 -331 321
rect -311 318 -307 321
rect -271 318 -267 321
rect -253 318 -249 321
rect -325 292 -321 298
rect -291 292 -287 298
rect -359 288 -333 292
rect -325 288 -299 292
rect -291 288 -277 292
rect -263 289 -259 298
rect -355 177 -351 288
rect -341 266 -338 288
rect -325 285 -321 288
rect -335 272 -331 275
rect -335 269 -321 272
rect -312 267 -289 271
rect -312 266 -308 267
rect -341 263 -308 266
rect -281 264 -277 288
rect -269 285 -259 289
rect -251 288 -243 292
rect -253 272 -249 275
rect -262 268 -249 272
rect -301 260 -258 264
rect -343 256 -309 260
rect -348 184 -344 255
rect -322 223 -319 256
rect -301 250 -297 260
rect -291 253 -267 257
rect -291 250 -287 253
rect -271 250 -267 253
rect -311 237 -307 240
rect -291 237 -287 240
rect -311 233 -287 237
rect -281 230 -277 240
rect -313 226 -266 230
rect -246 223 -243 288
rect -238 280 -235 319
rect -183 305 -163 309
rect -152 305 -94 309
rect -81 305 -61 309
rect -176 296 -172 305
rect -151 296 -147 305
rect -98 296 -94 305
rect -72 296 -68 305
rect -214 269 -173 273
rect -164 271 -160 289
rect -126 272 -122 289
rect -322 220 -243 223
rect -236 254 -194 258
rect -341 213 -287 217
rect -335 210 -331 213
rect -315 210 -311 213
rect -307 210 -303 213
rect -325 184 -321 190
rect -348 180 -333 184
rect -325 180 -311 184
rect -315 177 -311 180
rect -297 177 -293 190
rect -236 177 -232 254
rect -198 233 -194 254
rect -187 241 -183 269
rect -164 267 -136 271
rect -126 268 -109 272
rect -84 271 -80 289
rect -164 259 -160 267
rect -150 255 -122 259
rect -176 247 -172 250
rect -176 244 -165 247
rect -150 241 -146 255
rect -187 238 -146 241
rect -113 239 -109 268
rect -99 267 -80 271
rect -71 267 -59 271
rect -84 260 -80 267
rect -72 248 -68 251
rect -76 244 -68 248
rect -139 235 -98 239
rect -198 229 -148 233
rect -162 195 -158 229
rect -139 223 -135 235
rect -127 227 -95 232
rect -127 223 -122 227
rect -100 223 -95 227
rect -152 208 -147 213
rect -127 208 -122 213
rect -152 204 -122 208
rect -113 202 -109 213
rect -119 198 -109 202
rect -63 196 -59 267
rect -77 195 -59 196
rect -162 191 -59 195
rect -355 173 -323 177
rect -315 173 -305 177
rect -297 173 -232 177
rect -315 170 -311 173
rect -297 170 -293 173
rect -335 157 -331 160
rect -307 157 -303 160
rect -341 153 -287 157
rect -341 143 -243 147
rect -335 140 -331 143
rect -311 140 -307 143
rect -271 140 -267 143
rect -253 140 -249 143
rect -236 138 -232 173
rect -148 169 -110 174
rect -148 160 -143 169
rect -124 160 -120 169
rect -114 160 -110 169
rect -48 169 4 173
rect -133 140 -129 149
rect -236 137 -145 138
rect -236 135 -203 137
rect -198 135 -145 137
rect -133 136 -121 140
rect -102 136 -98 149
rect -48 159 -42 169
rect -1 159 4 169
rect -125 132 -110 136
rect -102 132 -43 136
rect -14 134 -9 148
rect -236 120 -224 121
rect -219 120 -132 121
rect -325 114 -321 120
rect -291 114 -287 120
rect -359 110 -333 114
rect -325 110 -299 114
rect -291 110 -277 114
rect -263 111 -259 120
rect -236 117 -132 120
rect -355 -1 -351 110
rect -341 88 -338 110
rect -325 107 -321 110
rect -335 94 -331 97
rect -335 91 -321 94
rect -312 89 -289 93
rect -312 88 -308 89
rect -341 85 -308 88
rect -281 86 -277 110
rect -269 107 -259 111
rect -251 110 -243 114
rect -253 94 -249 97
rect -262 90 -249 94
rect -301 82 -258 86
rect -343 78 -309 82
rect -348 6 -344 77
rect -322 45 -319 78
rect -301 72 -297 82
rect -291 75 -267 79
rect -291 72 -287 75
rect -271 72 -267 75
rect -311 59 -307 62
rect -291 59 -287 62
rect -311 55 -287 59
rect -281 52 -277 62
rect -313 48 -266 52
rect -246 45 -243 110
rect -236 87 -233 117
rect -125 108 -121 132
rect -102 109 -98 132
rect -14 129 3 134
rect -66 118 -25 122
rect -147 95 -143 100
rect -111 95 -107 101
rect -147 91 -107 95
rect -66 67 -62 118
rect -14 103 -9 129
rect -30 98 -9 103
rect 12 126 16 148
rect 56 139 76 143
rect 87 139 145 143
rect 158 139 178 143
rect 63 130 67 139
rect 88 130 92 139
rect 141 130 145 139
rect 167 130 171 139
rect 12 121 42 126
rect -30 95 -25 98
rect 12 95 16 121
rect 38 107 42 121
rect 38 103 66 107
rect 75 105 79 123
rect 113 106 117 123
rect -45 79 -40 87
rect -14 79 -9 87
rect 1 79 6 87
rect -45 74 6 79
rect 52 75 56 103
rect 75 101 103 105
rect 113 102 130 106
rect 155 105 159 123
rect 75 93 79 101
rect 89 89 117 93
rect 63 81 67 84
rect 63 78 74 81
rect 89 75 93 89
rect 52 72 93 75
rect 126 73 130 102
rect 140 101 159 105
rect 168 101 180 105
rect 155 94 159 101
rect 167 82 171 85
rect 163 78 171 82
rect 100 69 141 73
rect -322 42 -243 45
rect -233 62 -62 67
rect 53 63 91 67
rect -341 35 -287 39
rect -335 32 -331 35
rect -315 32 -311 35
rect -307 32 -303 35
rect -325 6 -321 12
rect -348 2 -333 6
rect -325 2 -311 6
rect -315 -1 -311 2
rect -297 -1 -293 12
rect -233 -1 -229 62
rect 53 46 57 63
rect -93 41 57 46
rect -203 -1 -199 32
rect -173 27 -135 32
rect -173 18 -168 27
rect -149 18 -145 27
rect -139 18 -135 27
rect 77 29 81 63
rect 100 57 104 69
rect 112 61 144 66
rect 112 57 117 61
rect 139 57 144 61
rect 87 42 92 47
rect 112 42 117 47
rect 87 38 117 42
rect 126 36 130 47
rect 120 32 130 36
rect 176 30 180 101
rect 162 29 180 30
rect 77 25 180 29
rect -355 -5 -323 -1
rect -315 -5 -305 -1
rect -297 -5 -229 -1
rect -315 -8 -311 -5
rect -297 -8 -293 -5
rect -335 -21 -331 -18
rect -307 -21 -303 -18
rect -341 -25 -282 -21
rect -233 -30 -229 -5
rect -215 -4 -199 -1
rect -158 -2 -154 7
rect -215 -5 -170 -4
rect -341 -35 -243 -31
rect -335 -38 -331 -35
rect -311 -38 -307 -35
rect -271 -38 -267 -35
rect -253 -38 -249 -35
rect -215 -46 -212 -5
rect -203 -8 -170 -5
rect -158 -6 -146 -2
rect -150 -10 -135 -6
rect -127 -8 -123 7
rect -90 13 -52 18
rect -90 4 -85 13
rect -66 4 -62 13
rect -56 4 -52 13
rect -173 -21 -160 -20
rect -173 -24 -157 -21
rect -162 -25 -157 -24
rect -150 -34 -146 -10
rect -127 -12 -105 -8
rect -127 -33 -123 -12
rect -108 -18 -105 -12
rect -75 -16 -71 -7
rect -108 -21 -87 -18
rect -75 -20 -63 -16
rect -67 -24 -52 -20
rect -44 -22 -40 -7
rect 11 -18 63 -14
rect -103 -39 -74 -36
rect -172 -47 -168 -42
rect -136 -47 -132 -41
rect -172 -51 -132 -47
rect -325 -64 -321 -58
rect -291 -64 -287 -58
rect -359 -68 -333 -64
rect -325 -68 -299 -64
rect -291 -68 -277 -64
rect -263 -67 -259 -58
rect -103 -59 -100 -39
rect -67 -48 -63 -24
rect -44 -26 -7 -22
rect -44 -47 -40 -26
rect -239 -62 -100 -59
rect -11 -50 -7 -26
rect 11 -28 17 -18
rect 58 -28 63 -18
rect 116 -22 136 -18
rect 147 -22 205 -18
rect 218 -22 238 -18
rect 123 -31 127 -22
rect 148 -31 152 -22
rect 201 -31 205 -22
rect 227 -31 231 -22
rect -11 -54 16 -50
rect 45 -53 50 -39
rect -89 -61 -85 -56
rect -53 -61 -49 -55
rect -355 -179 -351 -68
rect -341 -90 -338 -68
rect -325 -71 -321 -68
rect -335 -84 -331 -81
rect -335 -87 -321 -84
rect -312 -89 -289 -85
rect -312 -90 -308 -89
rect -341 -93 -308 -90
rect -281 -92 -277 -68
rect -269 -71 -259 -67
rect -251 -68 -243 -64
rect -253 -84 -249 -81
rect -262 -88 -249 -84
rect -301 -96 -258 -92
rect -343 -100 -309 -96
rect -348 -172 -344 -101
rect -322 -133 -319 -100
rect -301 -106 -297 -96
rect -291 -103 -267 -99
rect -291 -106 -287 -103
rect -271 -106 -267 -103
rect -311 -119 -307 -116
rect -291 -119 -287 -116
rect -311 -123 -287 -119
rect -281 -126 -277 -116
rect -313 -130 -266 -126
rect -246 -133 -243 -68
rect -239 -86 -235 -62
rect -89 -65 -49 -61
rect 45 -58 62 -53
rect -182 -71 -144 -66
rect -182 -80 -177 -71
rect -158 -80 -154 -71
rect -239 -89 -201 -86
rect -239 -91 -235 -89
rect -204 -119 -201 -89
rect -148 -80 -144 -71
rect 0 -68 34 -64
rect -167 -100 -163 -91
rect -189 -106 -179 -103
rect -167 -104 -155 -100
rect -159 -108 -144 -104
rect -136 -106 -132 -91
rect -90 -91 -38 -87
rect -90 -101 -84 -91
rect -43 -101 -38 -91
rect -204 -122 -166 -119
rect -322 -136 -243 -133
rect -237 -135 -226 -131
rect -159 -132 -155 -108
rect -136 -110 -104 -106
rect -136 -131 -132 -110
rect -107 -124 -104 -110
rect -107 -128 -85 -124
rect -56 -126 -51 -112
rect -341 -143 -287 -139
rect -335 -146 -331 -143
rect -315 -146 -311 -143
rect -307 -146 -303 -143
rect -237 -155 -233 -135
rect -56 -131 -39 -126
rect -30 -129 -26 -112
rect 0 -129 4 -68
rect 45 -84 50 -58
rect 29 -89 50 -84
rect 71 -60 75 -39
rect 97 -58 126 -54
rect 135 -56 139 -38
rect 173 -55 177 -38
rect 97 -60 101 -58
rect 71 -64 101 -60
rect 29 -92 34 -89
rect 71 -92 75 -64
rect 112 -86 116 -58
rect 135 -60 163 -56
rect 173 -59 190 -55
rect 215 -56 219 -38
rect 135 -68 139 -60
rect 149 -72 177 -68
rect 123 -80 127 -77
rect 123 -83 134 -80
rect 149 -86 153 -72
rect 112 -89 153 -86
rect 186 -88 190 -59
rect 200 -60 219 -56
rect 228 -60 240 -56
rect 215 -67 219 -60
rect 227 -79 231 -76
rect 223 -83 231 -79
rect 14 -108 19 -100
rect 45 -108 50 -100
rect 160 -92 201 -88
rect 137 -98 151 -94
rect 60 -108 65 -100
rect 14 -113 65 -108
rect -181 -145 -177 -140
rect -145 -145 -141 -139
rect -181 -149 -141 -145
rect -99 -142 -67 -138
rect -99 -161 -95 -142
rect -56 -157 -51 -131
rect -325 -172 -321 -166
rect -348 -176 -333 -172
rect -325 -176 -311 -172
rect -315 -179 -311 -176
rect -297 -179 -293 -166
rect -230 -163 -95 -161
rect -230 -164 -182 -163
rect -230 -179 -227 -164
rect -177 -164 -95 -163
rect -72 -162 -51 -157
rect -30 -133 4 -129
rect 137 -132 141 -98
rect 160 -104 164 -92
rect 172 -100 204 -95
rect 172 -104 177 -100
rect 199 -104 204 -100
rect 147 -119 152 -114
rect 172 -119 177 -114
rect 147 -123 177 -119
rect 186 -125 190 -114
rect 180 -129 190 -125
rect 236 -131 240 -60
rect 222 -132 240 -131
rect -72 -165 -67 -162
rect -30 -165 -26 -133
rect 137 -136 240 -132
rect 137 -148 140 -136
rect -355 -183 -323 -179
rect -315 -183 -305 -179
rect -297 -183 -227 -179
rect -87 -181 -82 -173
rect -56 -181 -51 -173
rect -9 -153 140 -148
rect -9 -163 -5 -153
rect -41 -181 -36 -173
rect -315 -186 -311 -183
rect -297 -186 -293 -183
rect -154 -190 -116 -185
rect -87 -186 -36 -181
rect -335 -199 -331 -196
rect -307 -199 -303 -196
rect -154 -199 -149 -190
rect -130 -199 -126 -190
rect -341 -203 -282 -199
rect -341 -213 -243 -209
rect -120 -199 -116 -190
rect -335 -216 -331 -213
rect -311 -216 -307 -213
rect -271 -216 -267 -213
rect -253 -216 -249 -213
rect -139 -219 -135 -210
rect -190 -224 -151 -221
rect -139 -223 -127 -219
rect -131 -227 -116 -223
rect -108 -225 -104 -210
rect -71 -204 -33 -199
rect -71 -213 -66 -204
rect -47 -213 -43 -204
rect -37 -213 -33 -204
rect 12 -212 50 -207
rect -325 -242 -321 -236
rect -291 -242 -287 -236
rect -359 -246 -333 -242
rect -325 -246 -299 -242
rect -291 -246 -277 -242
rect -263 -245 -259 -236
rect -211 -242 -138 -238
rect -355 -357 -351 -246
rect -341 -268 -338 -246
rect -325 -249 -321 -246
rect -335 -262 -331 -259
rect -335 -265 -321 -262
rect -312 -267 -289 -263
rect -312 -268 -308 -267
rect -341 -271 -308 -268
rect -281 -270 -277 -246
rect -269 -249 -259 -245
rect -251 -246 -243 -242
rect -253 -262 -249 -259
rect -262 -266 -249 -262
rect -301 -274 -258 -270
rect -343 -278 -309 -274
rect -348 -350 -344 -279
rect -322 -311 -319 -278
rect -301 -284 -297 -274
rect -291 -281 -267 -277
rect -291 -284 -287 -281
rect -271 -284 -267 -281
rect -311 -297 -307 -294
rect -291 -297 -287 -294
rect -311 -301 -287 -297
rect -281 -304 -277 -294
rect -313 -308 -266 -304
rect -246 -311 -243 -246
rect -131 -251 -127 -227
rect -108 -229 -86 -225
rect -108 -250 -104 -229
rect -89 -235 -86 -229
rect -56 -233 -52 -224
rect -89 -238 -68 -235
rect -56 -237 -44 -233
rect -48 -241 -33 -237
rect -25 -239 -21 -224
rect 12 -221 17 -212
rect 36 -221 40 -212
rect 46 -221 50 -212
rect -88 -255 -55 -252
rect -153 -264 -149 -259
rect -117 -264 -113 -258
rect -153 -268 -113 -264
rect -48 -265 -44 -241
rect -25 -243 -10 -239
rect 27 -241 31 -232
rect -25 -264 -21 -243
rect -13 -247 15 -243
rect 27 -245 39 -241
rect 35 -249 50 -245
rect 58 -247 62 -232
rect -233 -275 -229 -270
rect -232 -292 -229 -275
rect 3 -264 28 -260
rect -70 -278 -66 -273
rect -34 -278 -30 -272
rect -70 -282 -30 -278
rect 3 -292 6 -264
rect 35 -273 39 -249
rect 58 -251 73 -247
rect 58 -272 62 -251
rect 13 -286 17 -281
rect 49 -286 53 -280
rect 13 -290 53 -286
rect 69 -286 73 -251
rect 91 -254 143 -250
rect 91 -264 97 -254
rect 138 -264 143 -254
rect 69 -291 96 -286
rect 125 -289 130 -275
rect -232 -294 6 -292
rect -232 -296 -75 -294
rect -70 -296 6 -294
rect 125 -294 142 -289
rect -322 -314 -243 -311
rect -139 -306 -101 -301
rect -139 -315 -134 -306
rect -115 -315 -111 -306
rect -341 -321 -287 -317
rect -335 -324 -331 -321
rect -315 -324 -311 -321
rect -307 -324 -303 -321
rect -105 -315 -101 -306
rect 54 -305 114 -301
rect -325 -350 -321 -344
rect -348 -354 -333 -350
rect -325 -354 -311 -350
rect -315 -357 -311 -354
rect -297 -357 -293 -344
rect -124 -335 -120 -326
rect -228 -343 -223 -339
rect -164 -341 -136 -338
rect -124 -339 -112 -335
rect -164 -343 -161 -341
rect -228 -346 -161 -343
rect -116 -343 -101 -339
rect -93 -341 -89 -326
rect -56 -320 -18 -315
rect -56 -329 -51 -320
rect -32 -329 -28 -320
rect -22 -329 -18 -320
rect -355 -361 -323 -357
rect -315 -361 -305 -357
rect -297 -361 -228 -357
rect -196 -358 -123 -354
rect -315 -364 -311 -361
rect -297 -364 -293 -361
rect -335 -377 -331 -374
rect -307 -377 -303 -374
rect -341 -381 -282 -377
rect -232 -492 -228 -361
rect -116 -367 -112 -343
rect -93 -345 -71 -341
rect -93 -366 -89 -345
rect -74 -351 -71 -345
rect -41 -349 -37 -340
rect -10 -348 -6 -340
rect 54 -348 58 -305
rect 125 -320 130 -294
rect 109 -325 130 -320
rect 151 -321 155 -275
rect 151 -325 165 -321
rect 109 -328 114 -325
rect 151 -328 155 -325
rect -74 -354 -53 -351
rect -41 -353 -29 -349
rect -10 -352 58 -348
rect 94 -344 99 -336
rect 125 -344 130 -336
rect 140 -344 145 -336
rect 94 -349 145 -344
rect -33 -357 -18 -353
rect -65 -372 -40 -369
rect -138 -380 -134 -375
rect -102 -380 -98 -374
rect -138 -384 -98 -380
rect -33 -381 -29 -357
rect -10 -380 -6 -352
rect 161 -359 165 -325
rect 37 -363 165 -359
rect -55 -394 -51 -389
rect -19 -394 -15 -388
rect -141 -400 -103 -395
rect -55 -398 -15 -394
rect -141 -409 -136 -400
rect -117 -409 -113 -400
rect -107 -409 -103 -400
rect 37 -404 42 -363
rect 55 -371 107 -367
rect 55 -381 61 -371
rect 102 -381 107 -371
rect 37 -408 60 -404
rect 89 -406 94 -392
rect -126 -429 -122 -420
rect -173 -435 -138 -431
rect -126 -433 -114 -429
rect -118 -437 -103 -433
rect -95 -435 -91 -420
rect -46 -414 6 -410
rect -46 -424 -40 -414
rect 1 -424 6 -414
rect 89 -411 106 -406
rect 45 -422 78 -418
rect -212 -451 -125 -448
rect -118 -461 -114 -437
rect -95 -439 -67 -435
rect -95 -460 -91 -439
rect -71 -447 -67 -439
rect -71 -451 -41 -447
rect -12 -449 -7 -435
rect -12 -454 5 -449
rect -60 -465 -23 -460
rect -140 -474 -136 -469
rect -104 -474 -100 -468
rect -140 -478 -100 -474
rect -60 -492 -56 -465
rect -12 -480 -7 -454
rect -28 -485 -7 -480
rect 14 -459 18 -435
rect 45 -459 49 -422
rect 89 -437 94 -411
rect 73 -442 94 -437
rect 115 -419 119 -392
rect 115 -424 130 -419
rect 73 -445 78 -442
rect 115 -445 119 -424
rect 14 -464 49 -459
rect 58 -461 63 -453
rect 89 -461 94 -453
rect 104 -461 109 -453
rect -28 -488 -23 -485
rect 14 -488 18 -464
rect 58 -466 109 -461
rect -232 -497 -56 -492
rect -43 -504 -38 -496
rect -12 -504 -7 -496
rect 3 -504 8 -496
rect -43 -509 8 -504
<< m2contact >>
rect -348 255 -343 260
rect -258 259 -252 265
rect -240 275 -235 280
rect -219 268 -214 274
rect -98 235 -93 240
rect -203 132 -198 137
rect -224 120 -219 126
rect -348 77 -343 82
rect -258 81 -252 87
rect -236 82 -231 87
rect 141 69 146 74
rect -98 40 -93 46
rect -203 32 -198 39
rect -234 -36 -228 -30
rect -178 -24 -173 -19
rect -103 -36 -98 -31
rect -215 -51 -210 -46
rect -348 -101 -343 -96
rect -258 -97 -252 -91
rect -240 -96 -235 -91
rect -195 -106 -189 -101
rect -226 -135 -221 -130
rect 201 -92 206 -87
rect -238 -160 -233 -155
rect -182 -168 -177 -163
rect -9 -169 -4 -163
rect -195 -224 -190 -219
rect -216 -242 -211 -237
rect -348 -279 -343 -274
rect -258 -275 -252 -269
rect -93 -255 -88 -250
rect -238 -275 -233 -269
rect -9 -292 -4 -287
rect -217 -301 -212 -296
rect -75 -299 -70 -294
rect -228 -339 -223 -334
rect -201 -359 -196 -354
rect -70 -372 -65 -367
rect -218 -451 -212 -445
<< pdm12contact >>
rect -178 -435 -173 -430
<< metal2 >>
rect -362 256 -348 260
rect -240 264 -235 275
rect -252 260 -235 264
rect -224 126 -219 273
rect -54 239 -50 251
rect -93 235 -50 239
rect -359 78 -348 82
rect -252 82 -236 86
rect -241 -20 -237 82
rect -203 39 -198 132
rect 185 73 189 85
rect 146 69 189 73
rect -241 -23 -178 -20
rect -233 -39 -228 -36
rect -233 -42 -191 -39
rect -359 -100 -348 -96
rect -252 -96 -240 -92
rect -248 -147 -244 -96
rect -226 -130 -222 -42
rect -214 -133 -211 -51
rect -194 -101 -191 -42
rect -186 -54 -183 -23
rect -102 -31 -98 46
rect -186 -57 -104 -54
rect -214 -136 -192 -133
rect -248 -151 -212 -147
rect -238 -219 -234 -160
rect -238 -223 -224 -219
rect -359 -278 -348 -274
rect -252 -274 -238 -270
rect -228 -334 -224 -223
rect -216 -229 -212 -151
rect -195 -219 -192 -136
rect -216 -233 -197 -229
rect -216 -237 -212 -233
rect -217 -445 -213 -301
rect -201 -354 -197 -233
rect -182 -435 -178 -168
rect -107 -184 -104 -57
rect 245 -88 249 -76
rect 206 -92 249 -88
rect -107 -187 -90 -184
rect -93 -250 -90 -187
rect -9 -287 -5 -169
rect -74 -372 -70 -299
<< labels >>
rlabel metal1 -292 -308 -287 -304 1 gnd
rlabel metal1 -292 -130 -287 -126 1 gnd
rlabel metal1 -292 48 -287 52 1 gnd
rlabel metal1 -292 226 -287 230 1 gnd
rlabel metal1 -330 -265 -327 -262 1 gnd
rlabel metal1 -330 -87 -327 -84 1 gnd
rlabel metal1 -330 91 -327 94 1 gnd
rlabel metal1 -259 -265 -256 -262 1 gnd
rlabel metal1 -259 -87 -256 -84 1 gnd
rlabel metal1 -259 91 -256 94 1 gnd
rlabel metal1 -259 269 -256 272 1 gnd
rlabel metal1 -317 -213 -313 -209 4 vdd
rlabel metal1 -317 -35 -313 -31 4 vdd
rlabel metal1 -317 143 -313 147 4 vdd
rlabel metal1 -317 321 -313 325 4 vdd
rlabel metal1 -341 -321 -337 -317 4 vdd
rlabel metal1 -341 -143 -337 -139 4 vdd
rlabel metal1 -341 35 -337 39 4 vdd
rlabel metal1 -341 -381 -337 -377 2 gnd
rlabel metal1 -341 -203 -337 -199 2 gnd
rlabel metal1 -341 -25 -337 -21 2 gnd
rlabel metal1 -341 213 -337 217 4 vdd
rlabel metal1 -341 153 -337 157 2 gnd
rlabel metal1 -330 269 -326 272 1 gnd
rlabel metal1 -359 288 -355 292 3 a0
rlabel metal2 -362 256 -356 260 3 b0
rlabel metal1 -266 260 -262 264 1 p0
rlabel metal1 -284 173 -280 177 1 g0
rlabel metal1 -359 110 -356 114 3 a1
rlabel metal2 -359 78 -356 82 3 b1
rlabel metal2 -251 82 -247 86 1 p1
rlabel metal1 -282 -5 -276 -1 1 g1
rlabel metal2 -252 -96 -248 -92 1 p2
rlabel metal1 -359 -68 -356 -64 3 a2
rlabel metal2 -359 -100 -356 -96 3 b2
rlabel metal1 -359 -246 -356 -242 3 a3
rlabel metal1 -288 -183 -284 -179 1 g2
rlabel metal2 -359 -278 -356 -274 3 b3
rlabel metal2 -250 -274 -246 -270 1 p3
rlabel metal1 -287 -361 -283 -357 1 g3
rlabel metal1 -120 169 -114 174 5 vdd
rlabel metal1 -119 91 -114 95 1 gnd
rlabel metal1 -31 74 -25 79 1 gnd
rlabel metal1 -28 169 -17 173 5 vdd
rlabel metal1 16 121 20 126 1 c2
rlabel metal1 -61 -65 -56 -61 1 gnd
rlabel metal1 -62 13 -56 18 5 vdd
rlabel metal1 -144 -51 -139 -47 1 gnd
rlabel metal1 -145 27 -139 32 5 vdd
rlabel metal1 -154 -71 -148 -66 5 vdd
rlabel metal1 -153 -149 -148 -145 1 gnd
rlabel metal1 -70 -91 -59 -87 5 vdd
rlabel metal1 -73 -186 -67 -181 1 gnd
rlabel metal1 31 -18 42 -14 5 vdd
rlabel metal1 28 -113 34 -108 1 gnd
rlabel metal1 73 -64 78 -60 1 c3
rlabel metal1 -126 -190 -120 -185 5 vdd
rlabel metal1 -125 -268 -120 -264 1 gnd
rlabel metal1 -43 -204 -37 -199 5 vdd
rlabel metal1 -42 -282 -37 -278 1 gnd
rlabel metal1 40 -212 46 -207 5 vdd
rlabel metal1 41 -290 46 -286 1 gnd
rlabel metal1 -27 -398 -22 -394 1 gnd
rlabel metal1 -28 -320 -22 -315 5 vdd
rlabel metal1 -110 -384 -105 -380 1 gnd
rlabel metal1 -111 -306 -105 -301 5 vdd
rlabel metal1 -112 -478 -107 -474 1 gnd
rlabel metal1 -113 -400 -107 -395 5 vdd
rlabel metal1 111 -254 122 -250 5 vdd
rlabel metal1 108 -349 114 -344 1 gnd
rlabel metal1 75 -371 86 -367 5 vdd
rlabel metal1 72 -466 78 -461 1 gnd
rlabel metal1 -26 -414 -15 -410 5 vdd
rlabel metal1 -29 -509 -23 -504 1 gnd
rlabel metal1 122 -424 126 -419 1 c4
rlabel metal1 -168 305 -164 309 5 vdd
rlabel metal1 -119 198 -113 202 1 gnd
rlabel metal1 -76 244 -70 248 1 gnd
rlabel metal1 -176 244 -170 247 1 gnd
rlabel metal1 -76 305 -71 309 5 vdd
rlabel metal1 -139 305 -134 309 5 vdd
rlabel metal1 71 139 75 143 5 vdd
rlabel metal1 120 32 126 36 1 gnd
rlabel metal1 163 78 169 82 1 gnd
rlabel metal1 63 78 69 81 1 gnd
rlabel metal1 163 139 168 143 5 vdd
rlabel metal1 100 139 105 143 5 vdd
rlabel metal1 131 -22 135 -18 5 vdd
rlabel metal1 180 -129 186 -125 1 gnd
rlabel metal1 223 -83 229 -79 1 gnd
rlabel metal1 123 -83 129 -80 1 gnd
rlabel metal1 223 -22 228 -18 5 vdd
rlabel metal1 160 -22 165 -18 5 vdd
rlabel metal2 -54 245 -50 251 1 sum1
rlabel metal2 185 79 189 85 1 sum2
rlabel metal2 245 -82 249 -76 7 sum3
<< end >>
