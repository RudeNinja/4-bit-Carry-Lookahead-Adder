magic
tech scmos
timestamp 1638769712
<< nwell >>
rect 119 199 248 218
rect 139 55 201 78
<< ntransistor >>
rect 133 166 135 175
rect 225 167 227 176
rect 158 129 160 139
rect 170 129 172 139
rect 184 129 186 139
rect 197 129 199 139
rect 152 12 154 20
rect 165 12 167 20
rect 187 13 189 21
<< ptransistor >>
rect 133 205 135 212
rect 158 205 160 212
rect 170 205 172 212
rect 184 205 186 212
rect 197 205 199 212
rect 225 205 227 212
rect 152 61 154 72
rect 165 61 167 72
rect 187 61 189 72
<< ndiffusion >>
rect 130 166 133 175
rect 135 166 138 175
rect 222 167 225 176
rect 227 167 230 176
rect 155 129 158 139
rect 160 129 163 139
rect 167 129 170 139
rect 172 129 175 139
rect 180 129 184 139
rect 186 129 189 139
rect 193 129 197 139
rect 199 129 202 139
rect 207 129 209 139
rect 150 12 152 20
rect 154 12 165 20
rect 167 12 168 20
rect 186 13 187 21
rect 189 13 191 21
<< pdiffusion >>
rect 130 205 133 212
rect 135 205 138 212
rect 155 205 158 212
rect 160 205 170 212
rect 172 205 176 212
rect 180 205 184 212
rect 186 205 197 212
rect 199 205 204 212
rect 222 205 225 212
rect 227 205 230 212
rect 150 61 152 72
rect 154 61 160 72
rect 164 61 165 72
rect 167 61 169 72
rect 183 61 187 72
rect 189 61 191 72
<< ndcontact >>
rect 126 166 130 175
rect 138 166 142 175
rect 218 167 222 176
rect 230 167 234 176
rect 150 129 155 139
rect 163 129 167 139
rect 175 129 180 139
rect 189 129 193 139
rect 202 129 207 139
rect 146 12 150 20
rect 168 12 172 20
rect 182 13 186 21
rect 191 13 195 21
<< pdcontact >>
rect 126 205 130 212
rect 138 205 142 212
rect 151 205 155 212
rect 176 205 180 212
rect 204 205 208 212
rect 218 205 222 212
rect 230 205 234 212
rect 145 61 150 72
rect 160 61 164 72
rect 169 61 173 72
rect 179 61 183 72
rect 191 61 195 72
<< polysilicon >>
rect 133 212 135 215
rect 158 212 160 215
rect 170 212 172 215
rect 184 212 186 215
rect 197 212 199 215
rect 225 212 227 215
rect 133 175 135 205
rect 133 163 135 166
rect 158 139 160 205
rect 170 139 172 205
rect 184 139 186 205
rect 197 139 199 205
rect 225 176 227 205
rect 225 163 227 167
rect 158 126 160 129
rect 170 126 172 129
rect 184 126 186 129
rect 197 126 199 129
rect 152 72 154 75
rect 165 72 167 75
rect 187 72 189 75
rect 152 20 154 61
rect 165 20 167 61
rect 187 21 189 61
rect 152 9 154 12
rect 165 9 167 12
rect 187 10 189 13
<< polycontact >>
rect 129 185 133 189
rect 154 145 158 149
rect 166 183 170 187
rect 180 171 184 175
rect 199 183 203 187
rect 227 183 231 187
rect 148 46 152 50
rect 161 29 165 33
rect 183 44 187 48
<< metal1 >>
rect 119 221 139 225
rect 150 221 208 225
rect 221 221 241 225
rect 126 212 130 221
rect 151 212 155 221
rect 204 212 208 221
rect 230 212 234 221
rect 80 185 129 189
rect 138 187 142 205
rect 176 188 180 205
rect 83 33 87 185
rect 92 170 108 174
rect 95 50 99 170
rect 104 149 108 170
rect 115 157 119 185
rect 138 183 166 187
rect 176 184 193 188
rect 218 187 222 205
rect 138 175 142 183
rect 152 171 180 175
rect 126 163 130 166
rect 126 160 137 163
rect 152 157 156 171
rect 115 154 156 157
rect 189 155 193 184
rect 203 183 222 187
rect 231 183 243 187
rect 218 176 222 183
rect 230 164 234 167
rect 226 160 234 164
rect 163 151 204 155
rect 104 145 154 149
rect 140 111 144 145
rect 163 139 167 151
rect 175 143 207 148
rect 175 139 180 143
rect 202 139 207 143
rect 150 124 155 129
rect 175 124 180 129
rect 150 120 180 124
rect 189 118 193 129
rect 183 114 193 118
rect 239 112 243 183
rect 225 111 243 112
rect 140 107 243 111
rect 145 81 183 86
rect 145 72 150 81
rect 169 72 173 81
rect 179 72 183 81
rect 160 52 164 61
rect 95 46 148 50
rect 160 48 172 52
rect 168 44 183 48
rect 191 46 195 61
rect 83 29 161 33
rect 168 20 172 44
rect 191 42 203 46
rect 191 21 195 42
rect 146 7 150 12
rect 182 7 186 13
rect 146 3 186 7
<< m2contact >>
rect 204 151 209 156
<< metal2 >>
rect 248 155 252 165
rect 209 151 252 155
<< labels >>
rlabel metal1 134 221 138 225 5 vdd
rlabel metal1 183 114 189 118 1 gnd
rlabel metal1 226 160 232 164 1 gnd
rlabel metal1 126 160 132 163 1 gnd
rlabel metal1 226 221 231 225 5 vdd
rlabel metal1 163 221 168 225 5 vdd
rlabel metal1 173 81 179 86 5 vdd
rlabel metal1 174 3 179 7 1 gnd
rlabel metal2 248 160 252 165 1 propagate
rlabel metal1 199 42 203 46 1 generate
rlabel metal1 92 170 98 174 1 b
rlabel metal1 80 185 86 189 3 a
<< end >>
