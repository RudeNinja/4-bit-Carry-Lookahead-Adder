* SPICE3 file created from and_test2.ext - technology: scmos

.option scale=0.09u
.include TSMC_180nm.txt
.param SUPPLY=1.8

.global Gnd gnd vdd
Vdd vdd gnd 'SUPPLY'


vin_a1 a gnd pulse 0 1.8 0ns 100ps 100ps 9.9ns 20ns
vin_a2 b gnd pulse 0 1.8 0ns 100ps 100ps 19.9ns 40ns

M1000 a_n33_n13# a a_n45_n13# Gnd CMOSN w=8 l=2
+  ad=56 pd=30 as=80 ps=36
M1001 a_n45_n13# a vdd vdd CMOSP w=11 l=2
+  ad=77 pd=36 as=275 ps=116
M1002 gnd b a_n33_n13# Gnd CMOSN w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1003 out a_n45_n13# gnd Gnd CMOSN w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1004 vdd b a_n45_n13# vdd CMOSP w=11 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 out a_n45_n13# vdd vdd CMOSP w=11 l=2
+  ad=66 pd=34 as=0 ps=0
C0 vdd a 0.06fF
C1 a_n45_n13# vdd 0.16fF
C2 vdd b 0.06fF
C3 a_n45_n13# out 0.04fF
C4 a_n45_n13# a 0.08fF
C5 vdd vdd 0.11fF
C6 out gnd 0.07fF
C7 b a_n45_n13# 0.08fF
C8 b a 0.16fF
C9 vdd out 0.03fF
C10 vdd a_n45_n13# 0.09fF
C11 gnd Gnd 0.13fF
C12 out Gnd 0.16fF
C13 vdd Gnd 0.16fF
C14 a_n45_n13# Gnd 0.48fF
C15 b Gnd 0.25fF
C16 a Gnd 0.25fF
C17 vdd Gnd 1.43fF
.control
tran 0.1n 200n

set curplottitle= ShubhamPriyadarshan - 2020102027

plot v(a) v(b)+2 v(out)+4

.endc
.end