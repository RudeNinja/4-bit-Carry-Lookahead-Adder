magic
tech scmos
timestamp 1638820090
<< nwell >>
rect -804 731 -777 760
rect -559 722 -532 751
rect -298 746 -271 775
rect -894 635 -867 702
rect -789 635 -762 679
rect -894 583 -867 627
rect -789 583 -762 627
rect -649 626 -622 693
rect -544 626 -517 670
rect -388 650 -361 717
rect -283 650 -256 694
rect -649 574 -622 618
rect -544 574 -517 618
rect -388 598 -361 642
rect -283 598 -256 642
rect -209 521 -180 548
rect -128 536 -84 563
rect -76 536 -32 563
rect 80 536 124 563
rect 132 536 176 563
rect -894 427 -867 494
rect -789 427 -762 471
rect -894 375 -867 419
rect -789 375 -762 419
rect -649 418 -622 485
rect -544 418 -517 462
rect -388 442 -361 509
rect -283 442 -256 486
rect -649 366 -622 410
rect -544 366 -517 410
rect -388 390 -361 434
rect -283 390 -256 434
rect -151 431 -84 458
rect -76 431 -32 458
rect 57 431 124 458
rect 132 431 176 458
rect -922 284 -895 313
rect -831 261 -802 288
rect -750 276 -706 303
rect -698 276 -654 303
rect -542 276 -498 303
rect -490 276 -446 303
rect -341 292 -243 324
rect 65 316 94 343
rect 146 331 190 358
rect 198 331 242 358
rect 354 331 398 358
rect 406 331 450 358
rect -183 283 -54 302
rect -1012 188 -985 255
rect -907 188 -880 232
rect 123 226 190 253
rect 198 226 242 253
rect 331 226 398 253
rect 406 226 450 253
rect -1012 136 -985 180
rect -907 136 -880 180
rect -773 171 -706 198
rect -698 171 -654 198
rect -565 171 -498 198
rect -490 171 -446 198
rect -341 184 -287 216
rect -341 114 -243 146
rect -154 143 -92 166
rect -56 140 27 167
rect 56 117 185 136
rect 286 89 315 116
rect 367 104 411 131
rect 419 104 463 131
rect 575 104 619 131
rect 627 104 671 131
rect -844 47 -815 74
rect -763 62 -719 89
rect -711 62 -667 89
rect -555 62 -511 89
rect -503 62 -459 89
rect -1012 -20 -985 47
rect -907 -20 -880 24
rect -341 6 -287 38
rect -179 1 -117 24
rect -96 -13 -34 10
rect 344 -1 411 26
rect 419 -1 463 26
rect 552 -1 619 26
rect 627 -1 671 26
rect -1012 -72 -985 -28
rect -907 -72 -880 -28
rect -786 -43 -719 -16
rect -711 -43 -667 -16
rect -578 -43 -511 -16
rect -503 -43 -459 -16
rect -341 -64 -243 -32
rect 3 -47 86 -20
rect 116 -44 245 -25
rect -188 -97 -126 -74
rect -98 -120 -15 -93
rect 280 -125 309 -98
rect 361 -110 405 -83
rect 413 -110 457 -83
rect 569 -110 613 -83
rect 621 -110 665 -83
rect -846 -184 -817 -157
rect -765 -169 -721 -142
rect -713 -169 -669 -142
rect -557 -169 -513 -142
rect -505 -169 -461 -142
rect -341 -172 -287 -140
rect -341 -242 -243 -210
rect -160 -216 -98 -193
rect -77 -230 -15 -207
rect 338 -215 405 -188
rect 413 -215 457 -188
rect 546 -215 613 -188
rect 621 -215 665 -188
rect 6 -238 68 -215
rect -788 -274 -721 -247
rect -713 -274 -669 -247
rect -580 -274 -513 -247
rect -505 -274 -461 -247
rect 83 -283 166 -256
rect -341 -350 -287 -318
rect -145 -332 -83 -309
rect -62 -346 0 -323
rect 193 -349 222 -322
rect 274 -334 318 -307
rect 326 -334 370 -307
rect 482 -334 526 -307
rect 534 -334 578 -307
rect -855 -399 -826 -372
rect -774 -384 -730 -357
rect -722 -384 -678 -357
rect -566 -384 -522 -357
rect -514 -384 -470 -357
rect 47 -400 130 -373
rect -147 -426 -85 -403
rect -54 -443 29 -416
rect 251 -439 318 -412
rect 326 -439 370 -412
rect 459 -439 526 -412
rect 534 -439 578 -412
rect -797 -489 -730 -462
rect -722 -489 -678 -462
rect -589 -489 -522 -462
rect -514 -489 -470 -462
<< ntransistor >>
rect -325 760 -318 762
rect -831 745 -824 747
rect -586 736 -579 738
rect -415 702 -408 704
rect -921 687 -914 689
rect -676 678 -669 680
rect -440 677 -434 679
rect -335 677 -329 679
rect -946 662 -940 664
rect -841 662 -835 664
rect -440 662 -434 664
rect -335 662 -329 664
rect -701 653 -695 655
rect -596 653 -590 655
rect -946 647 -940 649
rect -841 647 -835 649
rect -701 638 -695 640
rect -596 638 -590 640
rect -440 625 -434 627
rect -335 625 -329 627
rect -946 610 -940 612
rect -841 610 -835 612
rect -440 610 -434 612
rect -335 610 -329 612
rect -701 601 -695 603
rect -596 601 -590 603
rect -946 595 -940 597
rect -841 595 -835 597
rect -701 586 -695 588
rect -596 586 -590 588
rect -415 494 -408 496
rect -196 494 -194 501
rect -113 484 -111 490
rect -98 484 -96 490
rect -61 484 -59 490
rect -46 484 -44 490
rect 95 484 97 490
rect 110 484 112 490
rect 147 484 149 490
rect 162 484 164 490
rect -921 479 -914 481
rect -676 470 -669 472
rect -440 469 -434 471
rect -335 469 -329 471
rect -946 454 -940 456
rect -841 454 -835 456
rect -440 454 -434 456
rect -335 454 -329 456
rect -701 445 -695 447
rect -596 445 -590 447
rect -946 439 -940 441
rect -841 439 -835 441
rect -701 430 -695 432
rect -596 430 -590 432
rect -440 417 -434 419
rect -335 417 -329 419
rect -138 404 -136 411
rect -946 402 -940 404
rect -841 402 -835 404
rect -440 402 -434 404
rect -335 402 -329 404
rect -701 393 -695 395
rect -596 393 -590 395
rect -946 387 -940 389
rect -841 387 -835 389
rect 70 404 72 411
rect -701 378 -695 380
rect -596 378 -590 380
rect -113 379 -111 385
rect -98 379 -96 385
rect -61 379 -59 385
rect -46 379 -44 385
rect 95 379 97 385
rect 110 379 112 385
rect 147 379 149 385
rect 162 379 164 385
rect -949 298 -942 300
rect -1039 240 -1032 242
rect -818 234 -816 241
rect -329 275 -327 285
rect 78 289 80 296
rect -257 275 -255 285
rect -169 250 -167 259
rect -305 240 -303 250
rect -295 240 -293 250
rect -285 240 -283 250
rect -275 240 -273 250
rect -735 224 -733 230
rect -720 224 -718 230
rect -683 224 -681 230
rect -668 224 -666 230
rect -527 224 -525 230
rect -512 224 -510 230
rect -475 224 -473 230
rect -460 224 -458 230
rect 161 279 163 285
rect 176 279 178 285
rect 213 279 215 285
rect 228 279 230 285
rect 369 279 371 285
rect 384 279 386 285
rect 421 279 423 285
rect 436 279 438 285
rect -77 251 -75 260
rect -1064 215 -1058 217
rect -959 215 -953 217
rect -144 213 -142 223
rect -132 213 -130 223
rect -118 213 -116 223
rect -105 213 -103 223
rect -1064 200 -1058 202
rect -959 200 -953 202
rect 136 199 138 206
rect -1064 163 -1058 165
rect -959 163 -953 165
rect -1064 148 -1058 150
rect -959 148 -953 150
rect -760 144 -758 151
rect -552 144 -550 151
rect 344 199 346 206
rect 161 174 163 180
rect 176 174 178 180
rect 213 174 215 180
rect 228 174 230 180
rect 369 174 371 180
rect 384 174 386 180
rect 421 174 423 180
rect 436 174 438 180
rect -329 160 -327 170
rect -319 160 -317 170
rect -301 160 -299 170
rect -735 119 -733 125
rect -720 119 -718 125
rect -683 119 -681 125
rect -668 119 -666 125
rect -527 119 -525 125
rect -512 119 -510 125
rect -475 119 -473 125
rect -460 119 -458 125
rect -329 97 -327 107
rect -257 97 -255 107
rect -141 100 -139 108
rect -128 100 -126 108
rect -106 101 -104 109
rect -38 87 -36 95
rect -20 87 -18 95
rect 7 87 9 95
rect 70 84 72 93
rect -1039 32 -1032 34
rect -831 20 -829 27
rect -305 62 -303 72
rect -295 62 -293 72
rect -285 62 -283 72
rect -275 62 -273 72
rect 162 85 164 94
rect 299 62 301 69
rect 95 47 97 57
rect 107 47 109 57
rect 121 47 123 57
rect 134 47 136 57
rect 382 52 384 58
rect 397 52 399 58
rect 434 52 436 58
rect 449 52 451 58
rect 590 52 592 58
rect 605 52 607 58
rect 642 52 644 58
rect 657 52 659 58
rect -748 10 -746 16
rect -733 10 -731 16
rect -696 10 -694 16
rect -681 10 -679 16
rect -540 10 -538 16
rect -525 10 -523 16
rect -488 10 -486 16
rect -473 10 -471 16
rect -1064 7 -1058 9
rect -959 7 -953 9
rect -1064 -8 -1058 -6
rect -959 -8 -953 -6
rect -329 -18 -327 -8
rect -319 -18 -317 -8
rect -301 -18 -299 -8
rect -1064 -45 -1058 -43
rect -959 -45 -953 -43
rect -1064 -60 -1058 -58
rect -959 -60 -953 -58
rect -773 -70 -771 -63
rect -565 -70 -563 -63
rect -166 -42 -164 -34
rect -153 -42 -151 -34
rect -131 -41 -129 -33
rect 357 -28 359 -21
rect -83 -56 -81 -48
rect -70 -56 -68 -48
rect -48 -55 -46 -47
rect -329 -81 -327 -71
rect -748 -95 -746 -89
rect -733 -95 -731 -89
rect -696 -95 -694 -89
rect -681 -95 -679 -89
rect -540 -95 -538 -89
rect -525 -95 -523 -89
rect -488 -95 -486 -89
rect -473 -95 -471 -89
rect -257 -81 -255 -71
rect -305 -116 -303 -106
rect -295 -116 -293 -106
rect -285 -116 -283 -106
rect -275 -116 -273 -106
rect 130 -77 132 -68
rect 21 -100 23 -92
rect 39 -100 41 -92
rect 66 -100 68 -92
rect 565 -28 567 -21
rect 382 -53 384 -47
rect 397 -53 399 -47
rect 434 -53 436 -47
rect 449 -53 451 -47
rect 590 -53 592 -47
rect 605 -53 607 -47
rect 642 -53 644 -47
rect 657 -53 659 -47
rect 222 -76 224 -67
rect -175 -140 -173 -132
rect -162 -140 -160 -132
rect -140 -139 -138 -131
rect -833 -211 -831 -204
rect 155 -114 157 -104
rect 167 -114 169 -104
rect 181 -114 183 -104
rect 194 -114 196 -104
rect 293 -152 295 -145
rect 376 -162 378 -156
rect 391 -162 393 -156
rect 428 -162 430 -156
rect 443 -162 445 -156
rect 584 -162 586 -156
rect 599 -162 601 -156
rect 636 -162 638 -156
rect 651 -162 653 -156
rect -80 -173 -78 -165
rect -62 -173 -60 -165
rect -35 -173 -33 -165
rect -329 -196 -327 -186
rect -319 -196 -317 -186
rect -301 -196 -299 -186
rect -750 -221 -748 -215
rect -735 -221 -733 -215
rect -698 -221 -696 -215
rect -683 -221 -681 -215
rect -542 -221 -540 -215
rect -527 -221 -525 -215
rect -490 -221 -488 -215
rect -475 -221 -473 -215
rect -329 -259 -327 -249
rect -775 -301 -773 -294
rect -567 -301 -565 -294
rect -257 -259 -255 -249
rect -147 -259 -145 -251
rect -134 -259 -132 -251
rect -112 -258 -110 -250
rect -64 -273 -62 -265
rect -51 -273 -49 -265
rect -29 -272 -27 -264
rect 351 -242 353 -235
rect 559 -242 561 -235
rect 19 -281 21 -273
rect 32 -281 34 -273
rect 54 -280 56 -272
rect 376 -267 378 -261
rect 391 -267 393 -261
rect 428 -267 430 -261
rect 443 -267 445 -261
rect 584 -267 586 -261
rect 599 -267 601 -261
rect 636 -267 638 -261
rect 651 -267 653 -261
rect -305 -294 -303 -284
rect -295 -294 -293 -284
rect -285 -294 -283 -284
rect -275 -294 -273 -284
rect -750 -326 -748 -320
rect -735 -326 -733 -320
rect -698 -326 -696 -320
rect -683 -326 -681 -320
rect -542 -326 -540 -320
rect -527 -326 -525 -320
rect -490 -326 -488 -320
rect -475 -326 -473 -320
rect -329 -374 -327 -364
rect -319 -374 -317 -364
rect -301 -374 -299 -364
rect 101 -336 103 -328
rect 119 -336 121 -328
rect 146 -336 148 -328
rect -132 -375 -130 -367
rect -119 -375 -117 -367
rect -97 -374 -95 -366
rect -842 -426 -840 -419
rect 206 -376 208 -369
rect -49 -389 -47 -381
rect -36 -389 -34 -381
rect -14 -388 -12 -380
rect 289 -386 291 -380
rect 304 -386 306 -380
rect 341 -386 343 -380
rect 356 -386 358 -380
rect 497 -386 499 -380
rect 512 -386 514 -380
rect 549 -386 551 -380
rect 564 -386 566 -380
rect -759 -436 -757 -430
rect -744 -436 -742 -430
rect -707 -436 -705 -430
rect -692 -436 -690 -430
rect -551 -436 -549 -430
rect -536 -436 -534 -430
rect -499 -436 -497 -430
rect -484 -436 -482 -430
rect -134 -469 -132 -461
rect -121 -469 -119 -461
rect -99 -468 -97 -460
rect -784 -516 -782 -509
rect -576 -516 -574 -509
rect 65 -453 67 -445
rect 83 -453 85 -445
rect 110 -453 112 -445
rect 264 -466 266 -459
rect 472 -466 474 -459
rect -36 -496 -34 -488
rect -18 -496 -16 -488
rect 9 -496 11 -488
rect 289 -491 291 -485
rect 304 -491 306 -485
rect 341 -491 343 -485
rect 356 -491 358 -485
rect 497 -491 499 -485
rect 512 -491 514 -485
rect 549 -491 551 -485
rect 564 -491 566 -485
rect -759 -541 -757 -535
rect -744 -541 -742 -535
rect -707 -541 -705 -535
rect -692 -541 -690 -535
rect -551 -541 -549 -535
rect -536 -541 -534 -535
rect -499 -541 -497 -535
rect -484 -541 -482 -535
<< ptransistor >>
rect -291 760 -279 762
rect -797 745 -785 747
rect -552 736 -540 738
rect -381 702 -369 704
rect -887 687 -875 689
rect -642 678 -630 680
rect -381 677 -369 679
rect -276 677 -264 679
rect -887 662 -875 664
rect -782 662 -770 664
rect -381 662 -369 664
rect -276 662 -264 664
rect -642 653 -630 655
rect -537 653 -525 655
rect -887 647 -875 649
rect -782 647 -770 649
rect -642 638 -630 640
rect -537 638 -525 640
rect -381 625 -369 627
rect -276 625 -264 627
rect -887 610 -875 612
rect -782 610 -770 612
rect -381 610 -369 612
rect -276 610 -264 612
rect -642 601 -630 603
rect -537 601 -525 603
rect -887 595 -875 597
rect -782 595 -770 597
rect -642 586 -630 588
rect -537 586 -525 588
rect -113 543 -111 555
rect -98 543 -96 555
rect -61 543 -59 555
rect -46 543 -44 555
rect 95 543 97 555
rect 110 543 112 555
rect 147 543 149 555
rect 162 543 164 555
rect -196 528 -194 540
rect -381 494 -369 496
rect -887 479 -875 481
rect -642 470 -630 472
rect -381 469 -369 471
rect -276 469 -264 471
rect -887 454 -875 456
rect -782 454 -770 456
rect -381 454 -369 456
rect -276 454 -264 456
rect -642 445 -630 447
rect -537 445 -525 447
rect -887 439 -875 441
rect -782 439 -770 441
rect -138 438 -136 450
rect -113 438 -111 450
rect -98 438 -96 450
rect -61 438 -59 450
rect -46 438 -44 450
rect 70 438 72 450
rect 95 438 97 450
rect 110 438 112 450
rect 147 438 149 450
rect 162 438 164 450
rect -642 430 -630 432
rect -537 430 -525 432
rect -381 417 -369 419
rect -276 417 -264 419
rect -887 402 -875 404
rect -782 402 -770 404
rect -381 402 -369 404
rect -276 402 -264 404
rect -642 393 -630 395
rect -537 393 -525 395
rect -887 387 -875 389
rect -782 387 -770 389
rect -642 378 -630 380
rect -537 378 -525 380
rect 161 338 163 350
rect 176 338 178 350
rect 213 338 215 350
rect 228 338 230 350
rect 369 338 371 350
rect 384 338 386 350
rect 421 338 423 350
rect 436 338 438 350
rect 78 323 80 335
rect -915 298 -903 300
rect -329 298 -327 318
rect -305 298 -303 318
rect -295 298 -293 318
rect -285 298 -283 318
rect -275 298 -273 318
rect -257 298 -255 318
rect -735 283 -733 295
rect -720 283 -718 295
rect -683 283 -681 295
rect -668 283 -666 295
rect -527 283 -525 295
rect -512 283 -510 295
rect -475 283 -473 295
rect -460 283 -458 295
rect -818 268 -816 280
rect -1005 240 -993 242
rect -169 289 -167 296
rect -144 289 -142 296
rect -132 289 -130 296
rect -118 289 -116 296
rect -105 289 -103 296
rect -77 289 -75 296
rect 136 233 138 245
rect 161 233 163 245
rect 176 233 178 245
rect 213 233 215 245
rect 228 233 230 245
rect 344 233 346 245
rect 369 233 371 245
rect 384 233 386 245
rect 421 233 423 245
rect 436 233 438 245
rect -1005 215 -993 217
rect -900 215 -888 217
rect -1005 200 -993 202
rect -900 200 -888 202
rect -329 190 -327 210
rect -319 190 -317 210
rect -301 190 -299 210
rect -760 178 -758 190
rect -735 178 -733 190
rect -720 178 -718 190
rect -683 178 -681 190
rect -668 178 -666 190
rect -552 178 -550 190
rect -527 178 -525 190
rect -512 178 -510 190
rect -475 178 -473 190
rect -460 178 -458 190
rect -1005 163 -993 165
rect -900 163 -888 165
rect -1005 148 -993 150
rect -900 148 -888 150
rect -141 149 -139 160
rect -128 149 -126 160
rect -106 149 -104 160
rect -329 120 -327 140
rect -305 120 -303 140
rect -295 120 -293 140
rect -285 120 -283 140
rect -275 120 -273 140
rect -257 120 -255 140
rect -748 69 -746 81
rect -733 69 -731 81
rect -696 69 -694 81
rect -681 69 -679 81
rect -540 69 -538 81
rect -525 69 -523 81
rect -488 69 -486 81
rect -473 69 -471 81
rect -38 148 -36 159
rect -20 148 -18 159
rect 7 148 9 159
rect 70 123 72 130
rect 95 123 97 130
rect 107 123 109 130
rect 121 123 123 130
rect 134 123 136 130
rect 162 123 164 130
rect -831 54 -829 66
rect -1005 32 -993 34
rect 382 111 384 123
rect 397 111 399 123
rect 434 111 436 123
rect 449 111 451 123
rect 590 111 592 123
rect 605 111 607 123
rect 642 111 644 123
rect 657 111 659 123
rect 299 96 301 108
rect -329 12 -327 32
rect -319 12 -317 32
rect -301 12 -299 32
rect -1005 7 -993 9
rect -900 7 -888 9
rect -1005 -8 -993 -6
rect -900 -8 -888 -6
rect -166 7 -164 18
rect -153 7 -151 18
rect -131 7 -129 18
rect -773 -36 -771 -24
rect -748 -36 -746 -24
rect -733 -36 -731 -24
rect -696 -36 -694 -24
rect -681 -36 -679 -24
rect -565 -36 -563 -24
rect -540 -36 -538 -24
rect -525 -36 -523 -24
rect -488 -36 -486 -24
rect -473 -36 -471 -24
rect 357 6 359 18
rect 382 6 384 18
rect 397 6 399 18
rect 434 6 436 18
rect 449 6 451 18
rect 565 6 567 18
rect 590 6 592 18
rect 605 6 607 18
rect 642 6 644 18
rect 657 6 659 18
rect -83 -7 -81 4
rect -70 -7 -68 4
rect -48 -7 -46 4
rect -1005 -45 -993 -43
rect -900 -45 -888 -43
rect -1005 -60 -993 -58
rect -900 -60 -888 -58
rect -329 -58 -327 -38
rect -305 -58 -303 -38
rect -295 -58 -293 -38
rect -285 -58 -283 -38
rect -275 -58 -273 -38
rect -257 -58 -255 -38
rect 21 -39 23 -28
rect 39 -39 41 -28
rect 66 -39 68 -28
rect 130 -38 132 -31
rect 155 -38 157 -31
rect 167 -38 169 -31
rect 181 -38 183 -31
rect 194 -38 196 -31
rect 222 -38 224 -31
rect -175 -91 -173 -80
rect -162 -91 -160 -80
rect -140 -91 -138 -80
rect -80 -112 -78 -101
rect -62 -112 -60 -101
rect -35 -112 -33 -101
rect 376 -103 378 -91
rect 391 -103 393 -91
rect 428 -103 430 -91
rect 443 -103 445 -91
rect 584 -103 586 -91
rect 599 -103 601 -91
rect 636 -103 638 -91
rect 651 -103 653 -91
rect -750 -162 -748 -150
rect -735 -162 -733 -150
rect -698 -162 -696 -150
rect -683 -162 -681 -150
rect -542 -162 -540 -150
rect -527 -162 -525 -150
rect -490 -162 -488 -150
rect -475 -162 -473 -150
rect -833 -177 -831 -165
rect -329 -166 -327 -146
rect -319 -166 -317 -146
rect -301 -166 -299 -146
rect 293 -118 295 -106
rect -147 -210 -145 -199
rect -134 -210 -132 -199
rect -112 -210 -110 -199
rect 351 -208 353 -196
rect 376 -208 378 -196
rect 391 -208 393 -196
rect 428 -208 430 -196
rect 443 -208 445 -196
rect 559 -208 561 -196
rect 584 -208 586 -196
rect 599 -208 601 -196
rect 636 -208 638 -196
rect 651 -208 653 -196
rect -329 -236 -327 -216
rect -305 -236 -303 -216
rect -295 -236 -293 -216
rect -285 -236 -283 -216
rect -275 -236 -273 -216
rect -257 -236 -255 -216
rect -775 -267 -773 -255
rect -750 -267 -748 -255
rect -735 -267 -733 -255
rect -698 -267 -696 -255
rect -683 -267 -681 -255
rect -567 -267 -565 -255
rect -542 -267 -540 -255
rect -527 -267 -525 -255
rect -490 -267 -488 -255
rect -475 -267 -473 -255
rect -64 -224 -62 -213
rect -51 -224 -49 -213
rect -29 -224 -27 -213
rect 19 -232 21 -221
rect 32 -232 34 -221
rect 54 -232 56 -221
rect 101 -275 103 -264
rect 119 -275 121 -264
rect 146 -275 148 -264
rect -329 -344 -327 -324
rect -319 -344 -317 -324
rect -301 -344 -299 -324
rect -132 -326 -130 -315
rect -119 -326 -117 -315
rect -97 -326 -95 -315
rect -759 -377 -757 -365
rect -744 -377 -742 -365
rect -707 -377 -705 -365
rect -692 -377 -690 -365
rect -551 -377 -549 -365
rect -536 -377 -534 -365
rect -499 -377 -497 -365
rect -484 -377 -482 -365
rect 289 -327 291 -315
rect 304 -327 306 -315
rect 341 -327 343 -315
rect 356 -327 358 -315
rect 497 -327 499 -315
rect 512 -327 514 -315
rect 549 -327 551 -315
rect 564 -327 566 -315
rect -49 -340 -47 -329
rect -36 -340 -34 -329
rect -14 -340 -12 -329
rect -842 -392 -840 -380
rect 206 -342 208 -330
rect 65 -392 67 -381
rect 83 -392 85 -381
rect 110 -392 112 -381
rect -134 -420 -132 -409
rect -121 -420 -119 -409
rect -99 -420 -97 -409
rect -36 -435 -34 -424
rect -18 -435 -16 -424
rect 9 -435 11 -424
rect -784 -482 -782 -470
rect -759 -482 -757 -470
rect -744 -482 -742 -470
rect -707 -482 -705 -470
rect -692 -482 -690 -470
rect -576 -482 -574 -470
rect -551 -482 -549 -470
rect -536 -482 -534 -470
rect -499 -482 -497 -470
rect -484 -482 -482 -470
rect 264 -432 266 -420
rect 289 -432 291 -420
rect 304 -432 306 -420
rect 341 -432 343 -420
rect 356 -432 358 -420
rect 472 -432 474 -420
rect 497 -432 499 -420
rect 512 -432 514 -420
rect 549 -432 551 -420
rect 564 -432 566 -420
<< ndiffusion >>
rect -325 762 -318 764
rect -325 756 -318 760
rect -831 747 -824 749
rect -831 741 -824 745
rect -586 738 -579 740
rect -586 732 -579 736
rect -415 704 -408 706
rect -415 698 -408 702
rect -921 689 -914 691
rect -921 683 -914 687
rect -676 680 -669 682
rect -440 679 -434 681
rect -335 679 -329 681
rect -676 674 -669 678
rect -946 664 -940 666
rect -841 664 -835 666
rect -440 664 -434 677
rect -335 664 -329 677
rect -946 649 -940 662
rect -841 649 -835 662
rect -701 655 -695 657
rect -596 655 -590 657
rect -440 659 -434 662
rect -335 659 -329 662
rect -946 644 -940 647
rect -841 644 -835 647
rect -701 640 -695 653
rect -596 640 -590 653
rect -701 635 -695 638
rect -596 635 -590 638
rect -440 627 -434 629
rect -335 627 -329 629
rect -946 612 -940 614
rect -841 612 -835 614
rect -440 612 -434 625
rect -335 612 -329 625
rect -946 597 -940 610
rect -841 597 -835 610
rect -701 603 -695 605
rect -596 603 -590 605
rect -440 607 -434 610
rect -335 607 -329 610
rect -946 592 -940 595
rect -841 592 -835 595
rect -701 588 -695 601
rect -596 588 -590 601
rect -701 583 -695 586
rect -596 583 -590 586
rect -415 496 -408 498
rect -198 494 -196 501
rect -194 494 -190 501
rect -415 490 -408 494
rect -921 481 -914 483
rect -115 484 -113 490
rect -111 484 -98 490
rect -96 484 -93 490
rect -63 484 -61 490
rect -59 484 -46 490
rect -44 484 -41 490
rect 93 484 95 490
rect 97 484 110 490
rect 112 484 115 490
rect 145 484 147 490
rect 149 484 162 490
rect 164 484 167 490
rect -921 475 -914 479
rect -676 472 -669 474
rect -440 471 -434 473
rect -335 471 -329 473
rect -676 466 -669 470
rect -946 456 -940 458
rect -841 456 -835 458
rect -440 456 -434 469
rect -335 456 -329 469
rect -946 441 -940 454
rect -841 441 -835 454
rect -701 447 -695 449
rect -596 447 -590 449
rect -440 451 -434 454
rect -335 451 -329 454
rect -946 436 -940 439
rect -841 436 -835 439
rect -701 432 -695 445
rect -596 432 -590 445
rect -701 427 -695 430
rect -596 427 -590 430
rect -440 419 -434 421
rect -335 419 -329 421
rect -946 404 -940 406
rect -841 404 -835 406
rect -440 404 -434 417
rect -335 404 -329 417
rect -140 404 -138 411
rect -136 404 -132 411
rect -946 389 -940 402
rect -841 389 -835 402
rect -701 395 -695 397
rect -596 395 -590 397
rect -440 399 -434 402
rect -335 399 -329 402
rect -946 384 -940 387
rect -841 384 -835 387
rect -701 380 -695 393
rect -596 380 -590 393
rect 68 404 70 411
rect 72 404 76 411
rect -115 379 -113 385
rect -111 379 -98 385
rect -96 379 -93 385
rect -63 379 -61 385
rect -59 379 -46 385
rect -44 379 -41 385
rect 93 379 95 385
rect 97 379 110 385
rect 112 379 115 385
rect 145 379 147 385
rect 149 379 162 385
rect 164 379 167 385
rect -701 375 -695 378
rect -596 375 -590 378
rect -949 300 -942 302
rect -949 294 -942 298
rect -1039 242 -1032 244
rect -1039 236 -1032 240
rect -820 234 -818 241
rect -816 234 -812 241
rect -331 275 -329 285
rect -327 275 -325 285
rect 76 289 78 296
rect 80 289 84 296
rect -259 275 -257 285
rect -255 275 -253 285
rect -172 250 -169 259
rect -167 250 -164 259
rect -307 240 -305 250
rect -303 240 -301 250
rect -297 240 -295 250
rect -293 240 -291 250
rect -287 240 -285 250
rect -283 240 -281 250
rect -277 240 -275 250
rect -273 240 -271 250
rect -737 224 -735 230
rect -733 224 -720 230
rect -718 224 -715 230
rect -685 224 -683 230
rect -681 224 -668 230
rect -666 224 -663 230
rect -529 224 -527 230
rect -525 224 -512 230
rect -510 224 -507 230
rect -477 224 -475 230
rect -473 224 -460 230
rect -458 224 -455 230
rect -1064 217 -1058 219
rect -959 217 -953 219
rect 159 279 161 285
rect 163 279 176 285
rect 178 279 181 285
rect 211 279 213 285
rect 215 279 228 285
rect 230 279 233 285
rect 367 279 369 285
rect 371 279 384 285
rect 386 279 389 285
rect 419 279 421 285
rect 423 279 436 285
rect 438 279 441 285
rect -80 251 -77 260
rect -75 251 -72 260
rect -1064 202 -1058 215
rect -959 202 -953 215
rect -147 213 -144 223
rect -142 213 -139 223
rect -135 213 -132 223
rect -130 213 -127 223
rect -122 213 -118 223
rect -116 213 -113 223
rect -109 213 -105 223
rect -103 213 -100 223
rect -95 213 -93 223
rect -1064 197 -1058 200
rect -959 197 -953 200
rect 134 199 136 206
rect 138 199 142 206
rect -1064 165 -1058 167
rect -959 165 -953 167
rect -1064 150 -1058 163
rect -959 150 -953 163
rect -1064 145 -1058 148
rect -959 145 -953 148
rect -762 144 -760 151
rect -758 144 -754 151
rect -554 144 -552 151
rect -550 144 -546 151
rect 342 199 344 206
rect 346 199 350 206
rect 159 174 161 180
rect 163 174 176 180
rect 178 174 181 180
rect 211 174 213 180
rect 215 174 228 180
rect 230 174 233 180
rect 367 174 369 180
rect 371 174 384 180
rect 386 174 389 180
rect 419 174 421 180
rect 423 174 436 180
rect 438 174 441 180
rect -331 160 -329 170
rect -327 160 -319 170
rect -317 160 -315 170
rect -303 160 -301 170
rect -299 160 -297 170
rect -737 119 -735 125
rect -733 119 -720 125
rect -718 119 -715 125
rect -685 119 -683 125
rect -681 119 -668 125
rect -666 119 -663 125
rect -529 119 -527 125
rect -525 119 -512 125
rect -510 119 -507 125
rect -477 119 -475 125
rect -473 119 -460 125
rect -458 119 -455 125
rect -331 97 -329 107
rect -327 97 -325 107
rect -259 97 -257 107
rect -255 97 -253 107
rect -143 100 -141 108
rect -139 100 -128 108
rect -126 100 -125 108
rect -107 101 -106 109
rect -104 101 -102 109
rect -40 87 -38 95
rect -36 87 -30 95
rect -25 87 -20 95
rect -18 87 -14 95
rect 6 87 7 95
rect 9 87 12 95
rect 67 84 70 93
rect 72 84 75 93
rect -1039 34 -1032 36
rect -1039 28 -1032 32
rect -833 20 -831 27
rect -829 20 -825 27
rect -307 62 -305 72
rect -303 62 -301 72
rect -297 62 -295 72
rect -293 62 -291 72
rect -287 62 -285 72
rect -283 62 -281 72
rect -277 62 -275 72
rect -273 62 -271 72
rect 159 85 162 94
rect 164 85 167 94
rect 297 62 299 69
rect 301 62 305 69
rect 92 47 95 57
rect 97 47 100 57
rect 104 47 107 57
rect 109 47 112 57
rect 117 47 121 57
rect 123 47 126 57
rect 130 47 134 57
rect 136 47 139 57
rect 144 47 146 57
rect 380 52 382 58
rect 384 52 397 58
rect 399 52 402 58
rect 432 52 434 58
rect 436 52 449 58
rect 451 52 454 58
rect 588 52 590 58
rect 592 52 605 58
rect 607 52 610 58
rect 640 52 642 58
rect 644 52 657 58
rect 659 52 662 58
rect -1064 9 -1058 11
rect -959 9 -953 11
rect -750 10 -748 16
rect -746 10 -733 16
rect -731 10 -728 16
rect -698 10 -696 16
rect -694 10 -681 16
rect -679 10 -676 16
rect -542 10 -540 16
rect -538 10 -525 16
rect -523 10 -520 16
rect -490 10 -488 16
rect -486 10 -473 16
rect -471 10 -468 16
rect -1064 -6 -1058 7
rect -959 -6 -953 7
rect -1064 -11 -1058 -8
rect -959 -11 -953 -8
rect -331 -18 -329 -8
rect -327 -18 -319 -8
rect -317 -18 -315 -8
rect -303 -18 -301 -8
rect -299 -18 -297 -8
rect -1064 -43 -1058 -41
rect -959 -43 -953 -41
rect -1064 -58 -1058 -45
rect -959 -58 -953 -45
rect -1064 -63 -1058 -60
rect -959 -63 -953 -60
rect -775 -70 -773 -63
rect -771 -70 -767 -63
rect -567 -70 -565 -63
rect -563 -70 -559 -63
rect -168 -42 -166 -34
rect -164 -42 -153 -34
rect -151 -42 -150 -34
rect -132 -41 -131 -33
rect -129 -41 -127 -33
rect 355 -28 357 -21
rect 359 -28 363 -21
rect -85 -56 -83 -48
rect -81 -56 -70 -48
rect -68 -56 -67 -48
rect -49 -55 -48 -47
rect -46 -55 -44 -47
rect -331 -81 -329 -71
rect -327 -81 -325 -71
rect -750 -95 -748 -89
rect -746 -95 -733 -89
rect -731 -95 -728 -89
rect -698 -95 -696 -89
rect -694 -95 -681 -89
rect -679 -95 -676 -89
rect -542 -95 -540 -89
rect -538 -95 -525 -89
rect -523 -95 -520 -89
rect -490 -95 -488 -89
rect -486 -95 -473 -89
rect -471 -95 -468 -89
rect -259 -81 -257 -71
rect -255 -81 -253 -71
rect -307 -116 -305 -106
rect -303 -116 -301 -106
rect -297 -116 -295 -106
rect -293 -116 -291 -106
rect -287 -116 -285 -106
rect -283 -116 -281 -106
rect -277 -116 -275 -106
rect -273 -116 -271 -106
rect 127 -77 130 -68
rect 132 -77 135 -68
rect 19 -100 21 -92
rect 23 -100 29 -92
rect 34 -100 39 -92
rect 41 -100 45 -92
rect 65 -100 66 -92
rect 68 -100 71 -92
rect 563 -28 565 -21
rect 567 -28 571 -21
rect 380 -53 382 -47
rect 384 -53 397 -47
rect 399 -53 402 -47
rect 432 -53 434 -47
rect 436 -53 449 -47
rect 451 -53 454 -47
rect 588 -53 590 -47
rect 592 -53 605 -47
rect 607 -53 610 -47
rect 640 -53 642 -47
rect 644 -53 657 -47
rect 659 -53 662 -47
rect 219 -76 222 -67
rect 224 -76 227 -67
rect -177 -140 -175 -132
rect -173 -140 -162 -132
rect -160 -140 -159 -132
rect -141 -139 -140 -131
rect -138 -139 -136 -131
rect -835 -211 -833 -204
rect -831 -211 -827 -204
rect 152 -114 155 -104
rect 157 -114 160 -104
rect 164 -114 167 -104
rect 169 -114 172 -104
rect 177 -114 181 -104
rect 183 -114 186 -104
rect 190 -114 194 -104
rect 196 -114 199 -104
rect 204 -114 206 -104
rect 291 -152 293 -145
rect 295 -152 299 -145
rect 374 -162 376 -156
rect 378 -162 391 -156
rect 393 -162 396 -156
rect 426 -162 428 -156
rect 430 -162 443 -156
rect 445 -162 448 -156
rect 582 -162 584 -156
rect 586 -162 599 -156
rect 601 -162 604 -156
rect 634 -162 636 -156
rect 638 -162 651 -156
rect 653 -162 656 -156
rect -82 -173 -80 -165
rect -78 -173 -72 -165
rect -67 -173 -62 -165
rect -60 -173 -56 -165
rect -36 -173 -35 -165
rect -33 -173 -30 -165
rect -331 -196 -329 -186
rect -327 -196 -319 -186
rect -317 -196 -315 -186
rect -303 -196 -301 -186
rect -299 -196 -297 -186
rect -752 -221 -750 -215
rect -748 -221 -735 -215
rect -733 -221 -730 -215
rect -700 -221 -698 -215
rect -696 -221 -683 -215
rect -681 -221 -678 -215
rect -544 -221 -542 -215
rect -540 -221 -527 -215
rect -525 -221 -522 -215
rect -492 -221 -490 -215
rect -488 -221 -475 -215
rect -473 -221 -470 -215
rect -331 -259 -329 -249
rect -327 -259 -325 -249
rect -777 -301 -775 -294
rect -773 -301 -769 -294
rect -569 -301 -567 -294
rect -565 -301 -561 -294
rect -259 -259 -257 -249
rect -255 -259 -253 -249
rect -149 -259 -147 -251
rect -145 -259 -134 -251
rect -132 -259 -131 -251
rect -113 -258 -112 -250
rect -110 -258 -108 -250
rect -66 -273 -64 -265
rect -62 -273 -51 -265
rect -49 -273 -48 -265
rect -30 -272 -29 -264
rect -27 -272 -25 -264
rect 349 -242 351 -235
rect 353 -242 357 -235
rect 557 -242 559 -235
rect 561 -242 565 -235
rect 17 -281 19 -273
rect 21 -281 32 -273
rect 34 -281 35 -273
rect 53 -280 54 -272
rect 56 -280 58 -272
rect 374 -267 376 -261
rect 378 -267 391 -261
rect 393 -267 396 -261
rect 426 -267 428 -261
rect 430 -267 443 -261
rect 445 -267 448 -261
rect 582 -267 584 -261
rect 586 -267 599 -261
rect 601 -267 604 -261
rect 634 -267 636 -261
rect 638 -267 651 -261
rect 653 -267 656 -261
rect -307 -294 -305 -284
rect -303 -294 -301 -284
rect -297 -294 -295 -284
rect -293 -294 -291 -284
rect -287 -294 -285 -284
rect -283 -294 -281 -284
rect -277 -294 -275 -284
rect -273 -294 -271 -284
rect -752 -326 -750 -320
rect -748 -326 -735 -320
rect -733 -326 -730 -320
rect -700 -326 -698 -320
rect -696 -326 -683 -320
rect -681 -326 -678 -320
rect -544 -326 -542 -320
rect -540 -326 -527 -320
rect -525 -326 -522 -320
rect -492 -326 -490 -320
rect -488 -326 -475 -320
rect -473 -326 -470 -320
rect -331 -374 -329 -364
rect -327 -374 -319 -364
rect -317 -374 -315 -364
rect -303 -374 -301 -364
rect -299 -374 -297 -364
rect 99 -336 101 -328
rect 103 -336 109 -328
rect 114 -336 119 -328
rect 121 -336 125 -328
rect 145 -336 146 -328
rect 148 -336 151 -328
rect -134 -375 -132 -367
rect -130 -375 -119 -367
rect -117 -375 -116 -367
rect -98 -374 -97 -366
rect -95 -374 -93 -366
rect -844 -426 -842 -419
rect -840 -426 -836 -419
rect 204 -376 206 -369
rect 208 -376 212 -369
rect -51 -389 -49 -381
rect -47 -389 -36 -381
rect -34 -389 -33 -381
rect -15 -388 -14 -380
rect -12 -388 -10 -380
rect 287 -386 289 -380
rect 291 -386 304 -380
rect 306 -386 309 -380
rect 339 -386 341 -380
rect 343 -386 356 -380
rect 358 -386 361 -380
rect 495 -386 497 -380
rect 499 -386 512 -380
rect 514 -386 517 -380
rect 547 -386 549 -380
rect 551 -386 564 -380
rect 566 -386 569 -380
rect -761 -436 -759 -430
rect -757 -436 -744 -430
rect -742 -436 -739 -430
rect -709 -436 -707 -430
rect -705 -436 -692 -430
rect -690 -436 -687 -430
rect -553 -436 -551 -430
rect -549 -436 -536 -430
rect -534 -436 -531 -430
rect -501 -436 -499 -430
rect -497 -436 -484 -430
rect -482 -436 -479 -430
rect -136 -469 -134 -461
rect -132 -469 -121 -461
rect -119 -469 -118 -461
rect -100 -468 -99 -460
rect -97 -468 -95 -460
rect -786 -516 -784 -509
rect -782 -516 -778 -509
rect -578 -516 -576 -509
rect -574 -516 -570 -509
rect 63 -453 65 -445
rect 67 -453 73 -445
rect 78 -453 83 -445
rect 85 -453 89 -445
rect 109 -453 110 -445
rect 112 -453 115 -445
rect 262 -466 264 -459
rect 266 -466 270 -459
rect 470 -466 472 -459
rect 474 -466 478 -459
rect -38 -496 -36 -488
rect -34 -496 -28 -488
rect -23 -496 -18 -488
rect -16 -496 -12 -488
rect 8 -496 9 -488
rect 11 -496 14 -488
rect 287 -491 289 -485
rect 291 -491 304 -485
rect 306 -491 309 -485
rect 339 -491 341 -485
rect 343 -491 356 -485
rect 358 -491 361 -485
rect 495 -491 497 -485
rect 499 -491 512 -485
rect 514 -491 517 -485
rect 547 -491 549 -485
rect 551 -491 564 -485
rect 566 -491 569 -485
rect -761 -541 -759 -535
rect -757 -541 -744 -535
rect -742 -541 -739 -535
rect -709 -541 -707 -535
rect -705 -541 -692 -535
rect -690 -541 -687 -535
rect -553 -541 -551 -535
rect -549 -541 -536 -535
rect -534 -541 -531 -535
rect -501 -541 -499 -535
rect -497 -541 -484 -535
rect -482 -541 -479 -535
<< pdiffusion >>
rect -291 762 -279 765
rect -291 756 -279 760
rect -797 747 -785 750
rect -797 741 -785 745
rect -552 738 -540 741
rect -552 732 -540 736
rect -381 704 -369 707
rect -381 698 -369 702
rect -887 689 -875 692
rect -887 683 -875 687
rect -642 680 -630 683
rect -381 679 -369 682
rect -276 679 -264 682
rect -887 664 -875 667
rect -642 674 -630 678
rect -782 664 -770 667
rect -381 673 -369 677
rect -381 664 -369 669
rect -276 673 -264 677
rect -276 664 -264 669
rect -887 658 -875 662
rect -887 649 -875 654
rect -782 658 -770 662
rect -642 655 -630 658
rect -537 655 -525 658
rect -381 660 -369 662
rect -276 660 -264 662
rect -782 649 -770 654
rect -887 645 -875 647
rect -782 645 -770 647
rect -642 649 -630 653
rect -642 640 -630 645
rect -537 649 -525 653
rect -537 640 -525 645
rect -642 636 -630 638
rect -537 636 -525 638
rect -381 627 -369 630
rect -276 627 -264 630
rect -887 612 -875 615
rect -782 612 -770 615
rect -381 621 -369 625
rect -381 612 -369 617
rect -276 621 -264 625
rect -276 612 -264 617
rect -887 606 -875 610
rect -887 597 -875 602
rect -782 606 -770 610
rect -642 603 -630 606
rect -537 603 -525 606
rect -381 608 -369 610
rect -276 608 -264 610
rect -782 597 -770 602
rect -887 593 -875 595
rect -782 593 -770 595
rect -642 597 -630 601
rect -642 588 -630 593
rect -537 597 -525 601
rect -537 588 -525 593
rect -642 584 -630 586
rect -537 584 -525 586
rect -116 543 -113 555
rect -111 543 -107 555
rect -103 543 -98 555
rect -96 543 -94 555
rect -64 543 -61 555
rect -59 543 -55 555
rect -51 543 -46 555
rect -44 543 -42 555
rect 92 543 95 555
rect 97 543 101 555
rect 105 543 110 555
rect 112 543 114 555
rect 144 543 147 555
rect 149 543 153 555
rect 157 543 162 555
rect 164 543 166 555
rect -199 528 -196 540
rect -194 528 -190 540
rect -381 496 -369 499
rect -381 490 -369 494
rect -887 481 -875 484
rect -887 475 -875 479
rect -642 472 -630 475
rect -381 471 -369 474
rect -276 471 -264 474
rect -887 456 -875 459
rect -642 466 -630 470
rect -782 456 -770 459
rect -381 465 -369 469
rect -381 456 -369 461
rect -276 465 -264 469
rect -276 456 -264 461
rect -887 450 -875 454
rect -887 441 -875 446
rect -782 450 -770 454
rect -642 447 -630 450
rect -537 447 -525 450
rect -381 452 -369 454
rect -276 452 -264 454
rect -782 441 -770 446
rect -887 437 -875 439
rect -782 437 -770 439
rect -642 441 -630 445
rect -642 432 -630 437
rect -537 441 -525 445
rect -141 438 -138 450
rect -136 438 -132 450
rect -116 438 -113 450
rect -111 438 -107 450
rect -103 438 -98 450
rect -96 438 -94 450
rect -64 438 -61 450
rect -59 438 -55 450
rect -51 438 -46 450
rect -44 438 -42 450
rect 67 438 70 450
rect 72 438 76 450
rect 92 438 95 450
rect 97 438 101 450
rect 105 438 110 450
rect 112 438 114 450
rect 144 438 147 450
rect 149 438 153 450
rect 157 438 162 450
rect 164 438 166 450
rect -537 432 -525 437
rect -642 428 -630 430
rect -537 428 -525 430
rect -381 419 -369 422
rect -276 419 -264 422
rect -887 404 -875 407
rect -782 404 -770 407
rect -381 413 -369 417
rect -381 404 -369 409
rect -276 413 -264 417
rect -276 404 -264 409
rect -887 398 -875 402
rect -887 389 -875 394
rect -782 398 -770 402
rect -642 395 -630 398
rect -537 395 -525 398
rect -381 400 -369 402
rect -276 400 -264 402
rect -782 389 -770 394
rect -887 385 -875 387
rect -782 385 -770 387
rect -642 389 -630 393
rect -642 380 -630 385
rect -537 389 -525 393
rect -537 380 -525 385
rect -642 376 -630 378
rect -537 376 -525 378
rect 158 338 161 350
rect 163 338 167 350
rect 171 338 176 350
rect 178 338 180 350
rect 210 338 213 350
rect 215 338 219 350
rect 223 338 228 350
rect 230 338 232 350
rect 366 338 369 350
rect 371 338 375 350
rect 379 338 384 350
rect 386 338 388 350
rect 418 338 421 350
rect 423 338 427 350
rect 431 338 436 350
rect 438 338 440 350
rect 75 323 78 335
rect 80 323 84 335
rect -915 300 -903 303
rect -331 298 -329 318
rect -327 298 -325 318
rect -307 298 -305 318
rect -303 298 -295 318
rect -293 298 -291 318
rect -287 298 -285 318
rect -283 298 -275 318
rect -273 298 -271 318
rect -259 298 -257 318
rect -255 298 -253 318
rect -915 294 -903 298
rect -738 283 -735 295
rect -733 283 -729 295
rect -725 283 -720 295
rect -718 283 -716 295
rect -686 283 -683 295
rect -681 283 -677 295
rect -673 283 -668 295
rect -666 283 -664 295
rect -530 283 -527 295
rect -525 283 -521 295
rect -517 283 -512 295
rect -510 283 -508 295
rect -478 283 -475 295
rect -473 283 -469 295
rect -465 283 -460 295
rect -458 283 -456 295
rect -821 268 -818 280
rect -816 268 -812 280
rect -1005 242 -993 245
rect -1005 236 -993 240
rect -172 289 -169 296
rect -167 289 -164 296
rect -147 289 -144 296
rect -142 289 -132 296
rect -130 289 -126 296
rect -122 289 -118 296
rect -116 289 -105 296
rect -103 289 -98 296
rect -80 289 -77 296
rect -75 289 -72 296
rect -1005 217 -993 220
rect 133 233 136 245
rect 138 233 142 245
rect 158 233 161 245
rect 163 233 167 245
rect 171 233 176 245
rect 178 233 180 245
rect 210 233 213 245
rect 215 233 219 245
rect 223 233 228 245
rect 230 233 232 245
rect 341 233 344 245
rect 346 233 350 245
rect 366 233 369 245
rect 371 233 375 245
rect 379 233 384 245
rect 386 233 388 245
rect 418 233 421 245
rect 423 233 427 245
rect 431 233 436 245
rect 438 233 440 245
rect -900 217 -888 220
rect -1005 211 -993 215
rect -1005 202 -993 207
rect -900 211 -888 215
rect -900 202 -888 207
rect -1005 198 -993 200
rect -900 198 -888 200
rect -331 190 -329 210
rect -327 190 -325 210
rect -321 190 -319 210
rect -317 190 -315 210
rect -303 190 -301 210
rect -299 190 -297 210
rect -763 178 -760 190
rect -758 178 -754 190
rect -738 178 -735 190
rect -733 178 -729 190
rect -725 178 -720 190
rect -718 178 -716 190
rect -686 178 -683 190
rect -681 178 -677 190
rect -673 178 -668 190
rect -666 178 -664 190
rect -555 178 -552 190
rect -550 178 -546 190
rect -530 178 -527 190
rect -525 178 -521 190
rect -517 178 -512 190
rect -510 178 -508 190
rect -478 178 -475 190
rect -473 178 -469 190
rect -465 178 -460 190
rect -458 178 -456 190
rect -1005 165 -993 168
rect -900 165 -888 168
rect -1005 159 -993 163
rect -1005 150 -993 155
rect -900 159 -888 163
rect -900 150 -888 155
rect -1005 146 -993 148
rect -900 146 -888 148
rect -143 149 -141 160
rect -139 149 -133 160
rect -129 149 -128 160
rect -126 149 -124 160
rect -110 149 -106 160
rect -104 149 -102 160
rect -331 120 -329 140
rect -327 120 -325 140
rect -307 120 -305 140
rect -303 120 -295 140
rect -293 120 -291 140
rect -287 120 -285 140
rect -283 120 -275 140
rect -273 120 -271 140
rect -259 120 -257 140
rect -255 120 -253 140
rect -751 69 -748 81
rect -746 69 -742 81
rect -738 69 -733 81
rect -731 69 -729 81
rect -699 69 -696 81
rect -694 69 -690 81
rect -686 69 -681 81
rect -679 69 -677 81
rect -543 69 -540 81
rect -538 69 -534 81
rect -530 69 -525 81
rect -523 69 -521 81
rect -491 69 -488 81
rect -486 69 -482 81
rect -478 69 -473 81
rect -471 69 -469 81
rect -42 148 -38 159
rect -36 148 -20 159
rect -18 148 -14 159
rect -4 148 -1 159
rect 4 148 7 159
rect 9 148 12 159
rect 16 148 18 159
rect 67 123 70 130
rect 72 123 75 130
rect 92 123 95 130
rect 97 123 107 130
rect 109 123 113 130
rect 117 123 121 130
rect 123 123 134 130
rect 136 123 141 130
rect 159 123 162 130
rect 164 123 167 130
rect -834 54 -831 66
rect -829 54 -825 66
rect -1005 34 -993 37
rect -1005 28 -993 32
rect 379 111 382 123
rect 384 111 388 123
rect 392 111 397 123
rect 399 111 401 123
rect 431 111 434 123
rect 436 111 440 123
rect 444 111 449 123
rect 451 111 453 123
rect 587 111 590 123
rect 592 111 596 123
rect 600 111 605 123
rect 607 111 609 123
rect 639 111 642 123
rect 644 111 648 123
rect 652 111 657 123
rect 659 111 661 123
rect 296 96 299 108
rect 301 96 305 108
rect -1005 9 -993 12
rect -900 9 -888 12
rect -331 12 -329 32
rect -327 12 -325 32
rect -321 12 -319 32
rect -317 12 -315 32
rect -303 12 -301 32
rect -299 12 -297 32
rect -1005 3 -993 7
rect -1005 -6 -993 -1
rect -900 3 -888 7
rect -900 -6 -888 -1
rect -168 7 -166 18
rect -164 7 -158 18
rect -154 7 -153 18
rect -151 7 -149 18
rect -135 7 -131 18
rect -129 7 -127 18
rect -1005 -10 -993 -8
rect -900 -10 -888 -8
rect -776 -36 -773 -24
rect -771 -36 -767 -24
rect -751 -36 -748 -24
rect -746 -36 -742 -24
rect -738 -36 -733 -24
rect -731 -36 -729 -24
rect -699 -36 -696 -24
rect -694 -36 -690 -24
rect -686 -36 -681 -24
rect -679 -36 -677 -24
rect -568 -36 -565 -24
rect -563 -36 -559 -24
rect -543 -36 -540 -24
rect -538 -36 -534 -24
rect -530 -36 -525 -24
rect -523 -36 -521 -24
rect -491 -36 -488 -24
rect -486 -36 -482 -24
rect -478 -36 -473 -24
rect -471 -36 -469 -24
rect 354 6 357 18
rect 359 6 363 18
rect 379 6 382 18
rect 384 6 388 18
rect 392 6 397 18
rect 399 6 401 18
rect 431 6 434 18
rect 436 6 440 18
rect 444 6 449 18
rect 451 6 453 18
rect 562 6 565 18
rect 567 6 571 18
rect 587 6 590 18
rect 592 6 596 18
rect 600 6 605 18
rect 607 6 609 18
rect 639 6 642 18
rect 644 6 648 18
rect 652 6 657 18
rect 659 6 661 18
rect -85 -7 -83 4
rect -81 -7 -75 4
rect -71 -7 -70 4
rect -68 -7 -66 4
rect -52 -7 -48 4
rect -46 -7 -44 4
rect -1005 -43 -993 -40
rect -900 -43 -888 -40
rect -1005 -49 -993 -45
rect -1005 -58 -993 -53
rect -900 -49 -888 -45
rect -900 -58 -888 -53
rect -1005 -62 -993 -60
rect -900 -62 -888 -60
rect -331 -58 -329 -38
rect -327 -58 -325 -38
rect -307 -58 -305 -38
rect -303 -58 -295 -38
rect -293 -58 -291 -38
rect -287 -58 -285 -38
rect -283 -58 -275 -38
rect -273 -58 -271 -38
rect -259 -58 -257 -38
rect -255 -58 -253 -38
rect 17 -39 21 -28
rect 23 -39 39 -28
rect 41 -39 45 -28
rect 55 -39 58 -28
rect 63 -39 66 -28
rect 68 -39 71 -28
rect 75 -39 77 -28
rect 127 -38 130 -31
rect 132 -38 135 -31
rect 152 -38 155 -31
rect 157 -38 167 -31
rect 169 -38 173 -31
rect 177 -38 181 -31
rect 183 -38 194 -31
rect 196 -38 201 -31
rect 219 -38 222 -31
rect 224 -38 227 -31
rect -177 -91 -175 -80
rect -173 -91 -167 -80
rect -163 -91 -162 -80
rect -160 -91 -158 -80
rect -144 -91 -140 -80
rect -138 -91 -136 -80
rect -84 -112 -80 -101
rect -78 -112 -62 -101
rect -60 -112 -56 -101
rect -46 -112 -43 -101
rect -38 -112 -35 -101
rect -33 -112 -30 -101
rect -26 -112 -24 -101
rect 373 -103 376 -91
rect 378 -103 382 -91
rect 386 -103 391 -91
rect 393 -103 395 -91
rect 425 -103 428 -91
rect 430 -103 434 -91
rect 438 -103 443 -91
rect 445 -103 447 -91
rect 581 -103 584 -91
rect 586 -103 590 -91
rect 594 -103 599 -91
rect 601 -103 603 -91
rect 633 -103 636 -91
rect 638 -103 642 -91
rect 646 -103 651 -91
rect 653 -103 655 -91
rect -753 -162 -750 -150
rect -748 -162 -744 -150
rect -740 -162 -735 -150
rect -733 -162 -731 -150
rect -701 -162 -698 -150
rect -696 -162 -692 -150
rect -688 -162 -683 -150
rect -681 -162 -679 -150
rect -545 -162 -542 -150
rect -540 -162 -536 -150
rect -532 -162 -527 -150
rect -525 -162 -523 -150
rect -493 -162 -490 -150
rect -488 -162 -484 -150
rect -480 -162 -475 -150
rect -473 -162 -471 -150
rect -836 -177 -833 -165
rect -831 -177 -827 -165
rect -331 -166 -329 -146
rect -327 -166 -325 -146
rect -321 -166 -319 -146
rect -317 -166 -315 -146
rect -303 -166 -301 -146
rect -299 -166 -297 -146
rect 290 -118 293 -106
rect 295 -118 299 -106
rect -149 -210 -147 -199
rect -145 -210 -139 -199
rect -135 -210 -134 -199
rect -132 -210 -130 -199
rect -116 -210 -112 -199
rect -110 -210 -108 -199
rect 348 -208 351 -196
rect 353 -208 357 -196
rect 373 -208 376 -196
rect 378 -208 382 -196
rect 386 -208 391 -196
rect 393 -208 395 -196
rect 425 -208 428 -196
rect 430 -208 434 -196
rect 438 -208 443 -196
rect 445 -208 447 -196
rect 556 -208 559 -196
rect 561 -208 565 -196
rect 581 -208 584 -196
rect 586 -208 590 -196
rect 594 -208 599 -196
rect 601 -208 603 -196
rect 633 -208 636 -196
rect 638 -208 642 -196
rect 646 -208 651 -196
rect 653 -208 655 -196
rect -331 -236 -329 -216
rect -327 -236 -325 -216
rect -307 -236 -305 -216
rect -303 -236 -295 -216
rect -293 -236 -291 -216
rect -287 -236 -285 -216
rect -283 -236 -275 -216
rect -273 -236 -271 -216
rect -259 -236 -257 -216
rect -255 -236 -253 -216
rect -778 -267 -775 -255
rect -773 -267 -769 -255
rect -753 -267 -750 -255
rect -748 -267 -744 -255
rect -740 -267 -735 -255
rect -733 -267 -731 -255
rect -701 -267 -698 -255
rect -696 -267 -692 -255
rect -688 -267 -683 -255
rect -681 -267 -679 -255
rect -570 -267 -567 -255
rect -565 -267 -561 -255
rect -545 -267 -542 -255
rect -540 -267 -536 -255
rect -532 -267 -527 -255
rect -525 -267 -523 -255
rect -493 -267 -490 -255
rect -488 -267 -484 -255
rect -480 -267 -475 -255
rect -473 -267 -471 -255
rect -66 -224 -64 -213
rect -62 -224 -56 -213
rect -52 -224 -51 -213
rect -49 -224 -47 -213
rect -33 -224 -29 -213
rect -27 -224 -25 -213
rect 17 -232 19 -221
rect 21 -232 27 -221
rect 31 -232 32 -221
rect 34 -232 36 -221
rect 50 -232 54 -221
rect 56 -232 58 -221
rect 97 -275 101 -264
rect 103 -275 119 -264
rect 121 -275 125 -264
rect 135 -275 138 -264
rect 143 -275 146 -264
rect 148 -275 151 -264
rect 155 -275 157 -264
rect -331 -344 -329 -324
rect -327 -344 -325 -324
rect -321 -344 -319 -324
rect -317 -344 -315 -324
rect -303 -344 -301 -324
rect -299 -344 -297 -324
rect -134 -326 -132 -315
rect -130 -326 -124 -315
rect -120 -326 -119 -315
rect -117 -326 -115 -315
rect -101 -326 -97 -315
rect -95 -326 -93 -315
rect -762 -377 -759 -365
rect -757 -377 -753 -365
rect -749 -377 -744 -365
rect -742 -377 -740 -365
rect -710 -377 -707 -365
rect -705 -377 -701 -365
rect -697 -377 -692 -365
rect -690 -377 -688 -365
rect -554 -377 -551 -365
rect -549 -377 -545 -365
rect -541 -377 -536 -365
rect -534 -377 -532 -365
rect -502 -377 -499 -365
rect -497 -377 -493 -365
rect -489 -377 -484 -365
rect -482 -377 -480 -365
rect 286 -327 289 -315
rect 291 -327 295 -315
rect 299 -327 304 -315
rect 306 -327 308 -315
rect 338 -327 341 -315
rect 343 -327 347 -315
rect 351 -327 356 -315
rect 358 -327 360 -315
rect 494 -327 497 -315
rect 499 -327 503 -315
rect 507 -327 512 -315
rect 514 -327 516 -315
rect 546 -327 549 -315
rect 551 -327 555 -315
rect 559 -327 564 -315
rect 566 -327 568 -315
rect -51 -340 -49 -329
rect -47 -340 -41 -329
rect -37 -340 -36 -329
rect -34 -340 -32 -329
rect -18 -340 -14 -329
rect -12 -340 -10 -329
rect -845 -392 -842 -380
rect -840 -392 -836 -380
rect 203 -342 206 -330
rect 208 -342 212 -330
rect 61 -392 65 -381
rect 67 -392 83 -381
rect 85 -392 89 -381
rect 99 -392 102 -381
rect 107 -392 110 -381
rect 112 -392 115 -381
rect 119 -392 121 -381
rect -136 -420 -134 -409
rect -132 -420 -126 -409
rect -122 -420 -121 -409
rect -119 -420 -117 -409
rect -103 -420 -99 -409
rect -97 -420 -95 -409
rect -40 -435 -36 -424
rect -34 -435 -18 -424
rect -16 -435 -12 -424
rect -2 -435 1 -424
rect 6 -435 9 -424
rect 11 -435 14 -424
rect 18 -435 20 -424
rect -787 -482 -784 -470
rect -782 -482 -778 -470
rect -762 -482 -759 -470
rect -757 -482 -753 -470
rect -749 -482 -744 -470
rect -742 -482 -740 -470
rect -710 -482 -707 -470
rect -705 -482 -701 -470
rect -697 -482 -692 -470
rect -690 -482 -688 -470
rect -579 -482 -576 -470
rect -574 -482 -570 -470
rect -554 -482 -551 -470
rect -549 -482 -545 -470
rect -541 -482 -536 -470
rect -534 -482 -532 -470
rect -502 -482 -499 -470
rect -497 -482 -493 -470
rect -489 -482 -484 -470
rect -482 -482 -480 -470
rect 261 -432 264 -420
rect 266 -432 270 -420
rect 286 -432 289 -420
rect 291 -432 295 -420
rect 299 -432 304 -420
rect 306 -432 308 -420
rect 338 -432 341 -420
rect 343 -432 347 -420
rect 351 -432 356 -420
rect 358 -432 360 -420
rect 469 -432 472 -420
rect 474 -432 478 -420
rect 494 -432 497 -420
rect 499 -432 503 -420
rect 507 -432 512 -420
rect 514 -432 516 -420
rect 546 -432 549 -420
rect 551 -432 555 -420
rect 559 -432 564 -420
rect 566 -432 568 -420
<< ndcontact >>
rect -325 764 -318 768
rect -831 749 -824 753
rect -325 752 -318 756
rect -831 737 -824 741
rect -586 740 -579 744
rect -586 728 -579 732
rect -415 706 -408 710
rect -921 691 -914 695
rect -415 694 -408 698
rect -921 679 -914 683
rect -676 682 -669 686
rect -440 681 -434 685
rect -335 681 -329 685
rect -946 666 -940 670
rect -841 666 -835 670
rect -676 670 -669 674
rect -701 657 -695 661
rect -596 657 -590 661
rect -440 655 -434 659
rect -335 655 -329 659
rect -946 640 -940 644
rect -841 640 -835 644
rect -701 631 -695 635
rect -596 631 -590 635
rect -440 629 -434 633
rect -335 629 -329 633
rect -946 614 -940 618
rect -841 614 -835 618
rect -701 605 -695 609
rect -596 605 -590 609
rect -440 603 -434 607
rect -335 603 -329 607
rect -946 588 -940 592
rect -841 588 -835 592
rect -701 579 -695 583
rect -596 579 -590 583
rect -415 498 -408 502
rect -202 494 -198 501
rect -190 494 -186 501
rect -921 483 -914 487
rect -415 486 -408 490
rect -119 484 -115 490
rect -93 484 -89 490
rect -67 484 -63 490
rect -41 484 -37 490
rect 89 484 93 490
rect 115 484 119 490
rect 141 484 145 490
rect 167 484 171 490
rect -921 471 -914 475
rect -676 474 -669 478
rect -440 473 -434 477
rect -335 473 -329 477
rect -946 458 -940 462
rect -841 458 -835 462
rect -676 462 -669 466
rect -701 449 -695 453
rect -596 449 -590 453
rect -440 447 -434 451
rect -335 447 -329 451
rect -946 432 -940 436
rect -841 432 -835 436
rect -701 423 -695 427
rect -596 423 -590 427
rect -440 421 -434 425
rect -335 421 -329 425
rect -946 406 -940 410
rect -841 406 -835 410
rect -144 404 -140 411
rect -132 404 -128 411
rect -701 397 -695 401
rect -596 397 -590 401
rect -440 395 -434 399
rect -335 395 -329 399
rect -946 380 -940 384
rect -841 380 -835 384
rect 64 404 68 411
rect 76 404 80 411
rect -119 379 -115 385
rect -93 379 -89 385
rect -67 379 -63 385
rect -41 379 -37 385
rect 89 379 93 385
rect 115 379 119 385
rect 141 379 145 385
rect 167 379 171 385
rect -701 371 -695 375
rect -596 371 -590 375
rect -949 302 -942 306
rect -949 290 -942 294
rect -1039 244 -1032 248
rect -1039 232 -1032 236
rect -824 234 -820 241
rect -812 234 -808 241
rect -335 275 -331 285
rect -325 275 -321 285
rect 72 289 76 296
rect 84 289 88 296
rect -263 275 -259 285
rect -253 275 -249 285
rect -176 250 -172 259
rect -164 250 -160 259
rect -311 240 -307 250
rect -301 240 -297 250
rect -291 240 -287 250
rect -281 240 -277 250
rect -271 240 -267 250
rect -741 224 -737 230
rect -715 224 -711 230
rect -689 224 -685 230
rect -663 224 -659 230
rect -533 224 -529 230
rect -507 224 -503 230
rect -481 224 -477 230
rect -455 224 -451 230
rect -1064 219 -1058 223
rect -959 219 -953 223
rect 155 279 159 285
rect 181 279 185 285
rect 207 279 211 285
rect 233 279 237 285
rect 363 279 367 285
rect 389 279 393 285
rect 415 279 419 285
rect 441 279 445 285
rect -84 251 -80 260
rect -72 251 -68 260
rect -152 213 -147 223
rect -139 213 -135 223
rect -127 213 -122 223
rect -113 213 -109 223
rect -100 213 -95 223
rect -1064 193 -1058 197
rect -959 193 -953 197
rect 130 199 134 206
rect 142 199 146 206
rect -1064 167 -1058 171
rect -959 167 -953 171
rect -1064 141 -1058 145
rect -959 141 -953 145
rect -766 144 -762 151
rect -754 144 -750 151
rect -558 144 -554 151
rect -546 144 -542 151
rect 338 199 342 206
rect 350 199 354 206
rect 155 174 159 180
rect 181 174 185 180
rect 207 174 211 180
rect 233 174 237 180
rect 363 174 367 180
rect 389 174 393 180
rect 415 174 419 180
rect 441 174 445 180
rect -335 160 -331 170
rect -315 160 -311 170
rect -307 160 -303 170
rect -297 160 -293 170
rect -741 119 -737 125
rect -715 119 -711 125
rect -689 119 -685 125
rect -663 119 -659 125
rect -533 119 -529 125
rect -507 119 -503 125
rect -481 119 -477 125
rect -455 119 -451 125
rect -335 97 -331 107
rect -325 97 -321 107
rect -263 97 -259 107
rect -253 97 -249 107
rect -147 100 -143 108
rect -125 100 -121 108
rect -111 101 -107 109
rect -102 101 -98 109
rect -45 87 -40 95
rect -30 87 -25 95
rect -14 87 -9 95
rect 1 87 6 95
rect 12 87 16 95
rect 63 84 67 93
rect 75 84 79 93
rect -1039 36 -1032 40
rect -1039 24 -1032 28
rect -837 20 -833 27
rect -825 20 -821 27
rect -311 62 -307 72
rect -301 62 -297 72
rect -291 62 -287 72
rect -281 62 -277 72
rect -271 62 -267 72
rect 155 85 159 94
rect 167 85 171 94
rect 293 62 297 69
rect 305 62 309 69
rect 87 47 92 57
rect 100 47 104 57
rect 112 47 117 57
rect 126 47 130 57
rect 139 47 144 57
rect 376 52 380 58
rect 402 52 406 58
rect 428 52 432 58
rect 454 52 458 58
rect 584 52 588 58
rect 610 52 614 58
rect 636 52 640 58
rect 662 52 666 58
rect -1064 11 -1058 15
rect -959 11 -953 15
rect -754 10 -750 16
rect -728 10 -724 16
rect -702 10 -698 16
rect -676 10 -672 16
rect -546 10 -542 16
rect -520 10 -516 16
rect -494 10 -490 16
rect -468 10 -464 16
rect -1064 -15 -1058 -11
rect -959 -15 -953 -11
rect -335 -18 -331 -8
rect -315 -18 -311 -8
rect -307 -18 -303 -8
rect -297 -18 -293 -8
rect -1064 -41 -1058 -37
rect -959 -41 -953 -37
rect -1064 -67 -1058 -63
rect -959 -67 -953 -63
rect -779 -70 -775 -63
rect -767 -70 -763 -63
rect -571 -70 -567 -63
rect -559 -70 -555 -63
rect -172 -42 -168 -34
rect -150 -42 -146 -34
rect -136 -41 -132 -33
rect -127 -41 -123 -33
rect 351 -28 355 -21
rect 363 -28 367 -21
rect -89 -56 -85 -48
rect -67 -56 -63 -48
rect -53 -55 -49 -47
rect -44 -55 -40 -47
rect -335 -81 -331 -71
rect -325 -81 -321 -71
rect -754 -95 -750 -89
rect -728 -95 -724 -89
rect -702 -95 -698 -89
rect -676 -95 -672 -89
rect -546 -95 -542 -89
rect -520 -95 -516 -89
rect -494 -95 -490 -89
rect -468 -95 -464 -89
rect -263 -81 -259 -71
rect -253 -81 -249 -71
rect -311 -116 -307 -106
rect -301 -116 -297 -106
rect -291 -116 -287 -106
rect -281 -116 -277 -106
rect -271 -116 -267 -106
rect 123 -77 127 -68
rect 135 -77 139 -68
rect 14 -100 19 -92
rect 29 -100 34 -92
rect 45 -100 50 -92
rect 60 -100 65 -92
rect 71 -100 75 -92
rect 559 -28 563 -21
rect 571 -28 575 -21
rect 376 -53 380 -47
rect 402 -53 406 -47
rect 428 -53 432 -47
rect 454 -53 458 -47
rect 584 -53 588 -47
rect 610 -53 614 -47
rect 636 -53 640 -47
rect 662 -53 666 -47
rect 215 -76 219 -67
rect 227 -76 231 -67
rect -181 -140 -177 -132
rect -159 -140 -155 -132
rect -145 -139 -141 -131
rect -136 -139 -132 -131
rect -839 -211 -835 -204
rect -827 -211 -823 -204
rect 147 -114 152 -104
rect 160 -114 164 -104
rect 172 -114 177 -104
rect 186 -114 190 -104
rect 199 -114 204 -104
rect 287 -152 291 -145
rect 299 -152 303 -145
rect 370 -162 374 -156
rect 396 -162 400 -156
rect 422 -162 426 -156
rect 448 -162 452 -156
rect 578 -162 582 -156
rect 604 -162 608 -156
rect 630 -162 634 -156
rect 656 -162 660 -156
rect -87 -173 -82 -165
rect -72 -173 -67 -165
rect -56 -173 -51 -165
rect -41 -173 -36 -165
rect -30 -173 -26 -165
rect -335 -196 -331 -186
rect -315 -196 -311 -186
rect -307 -196 -303 -186
rect -297 -196 -293 -186
rect -756 -221 -752 -215
rect -730 -221 -726 -215
rect -704 -221 -700 -215
rect -678 -221 -674 -215
rect -548 -221 -544 -215
rect -522 -221 -518 -215
rect -496 -221 -492 -215
rect -470 -221 -466 -215
rect -335 -259 -331 -249
rect -325 -259 -321 -249
rect -781 -301 -777 -294
rect -769 -301 -765 -294
rect -573 -301 -569 -294
rect -561 -301 -557 -294
rect -263 -259 -259 -249
rect -253 -259 -249 -249
rect -153 -259 -149 -251
rect -131 -259 -127 -251
rect -117 -258 -113 -250
rect -108 -258 -104 -250
rect -70 -273 -66 -265
rect -48 -273 -44 -265
rect -34 -272 -30 -264
rect -25 -272 -21 -264
rect 345 -242 349 -235
rect 357 -242 361 -235
rect 553 -242 557 -235
rect 565 -242 569 -235
rect 13 -281 17 -273
rect 35 -281 39 -273
rect 49 -280 53 -272
rect 58 -280 62 -272
rect 370 -267 374 -261
rect 396 -267 400 -261
rect 422 -267 426 -261
rect 448 -267 452 -261
rect 578 -267 582 -261
rect 604 -267 608 -261
rect 630 -267 634 -261
rect 656 -267 660 -261
rect -311 -294 -307 -284
rect -301 -294 -297 -284
rect -291 -294 -287 -284
rect -281 -294 -277 -284
rect -271 -294 -267 -284
rect -756 -326 -752 -320
rect -730 -326 -726 -320
rect -704 -326 -700 -320
rect -678 -326 -674 -320
rect -548 -326 -544 -320
rect -522 -326 -518 -320
rect -496 -326 -492 -320
rect -470 -326 -466 -320
rect -335 -374 -331 -364
rect -315 -374 -311 -364
rect -307 -374 -303 -364
rect -297 -374 -293 -364
rect 94 -336 99 -328
rect 109 -336 114 -328
rect 125 -336 130 -328
rect 140 -336 145 -328
rect 151 -336 155 -328
rect -138 -375 -134 -367
rect -116 -375 -112 -367
rect -102 -374 -98 -366
rect -93 -374 -89 -366
rect -848 -426 -844 -419
rect -836 -426 -832 -419
rect 200 -376 204 -369
rect 212 -376 216 -369
rect -55 -389 -51 -381
rect -33 -389 -29 -381
rect -19 -388 -15 -380
rect -10 -388 -6 -380
rect 283 -386 287 -380
rect 309 -386 313 -380
rect 335 -386 339 -380
rect 361 -386 365 -380
rect 491 -386 495 -380
rect 517 -386 521 -380
rect 543 -386 547 -380
rect 569 -386 573 -380
rect -765 -436 -761 -430
rect -739 -436 -735 -430
rect -713 -436 -709 -430
rect -687 -436 -683 -430
rect -557 -436 -553 -430
rect -531 -436 -527 -430
rect -505 -436 -501 -430
rect -479 -436 -475 -430
rect -140 -469 -136 -461
rect -118 -469 -114 -461
rect -104 -468 -100 -460
rect -95 -468 -91 -460
rect -790 -516 -786 -509
rect -778 -516 -774 -509
rect -582 -516 -578 -509
rect -570 -516 -566 -509
rect 58 -453 63 -445
rect 73 -453 78 -445
rect 89 -453 94 -445
rect 104 -453 109 -445
rect 115 -453 119 -445
rect 258 -466 262 -459
rect 270 -466 274 -459
rect 466 -466 470 -459
rect 478 -466 482 -459
rect -43 -496 -38 -488
rect -28 -496 -23 -488
rect -12 -496 -7 -488
rect 3 -496 8 -488
rect 14 -496 18 -488
rect 283 -491 287 -485
rect 309 -491 313 -485
rect 335 -491 339 -485
rect 361 -491 365 -485
rect 491 -491 495 -485
rect 517 -491 521 -485
rect 543 -491 547 -485
rect 569 -491 573 -485
rect -765 -541 -761 -535
rect -739 -541 -735 -535
rect -713 -541 -709 -535
rect -687 -541 -683 -535
rect -557 -541 -553 -535
rect -531 -541 -527 -535
rect -505 -541 -501 -535
rect -479 -541 -475 -535
<< pdcontact >>
rect -291 765 -279 769
rect -797 750 -785 754
rect -291 752 -279 756
rect -797 737 -785 741
rect -552 741 -540 745
rect -552 728 -540 732
rect -381 707 -369 711
rect -887 692 -875 696
rect -381 694 -369 698
rect -887 679 -875 683
rect -642 683 -630 687
rect -381 682 -369 686
rect -276 682 -264 686
rect -887 667 -875 671
rect -782 667 -770 671
rect -642 670 -630 674
rect -381 669 -369 673
rect -276 669 -264 673
rect -887 654 -875 658
rect -782 654 -770 658
rect -642 658 -630 662
rect -537 658 -525 662
rect -381 656 -369 660
rect -276 656 -264 660
rect -887 641 -875 645
rect -782 641 -770 645
rect -642 645 -630 649
rect -537 645 -525 649
rect -642 632 -630 636
rect -537 632 -525 636
rect -381 630 -369 634
rect -276 630 -264 634
rect -887 615 -875 619
rect -782 615 -770 619
rect -381 617 -369 621
rect -276 617 -264 621
rect -887 602 -875 606
rect -782 602 -770 606
rect -642 606 -630 610
rect -537 606 -525 610
rect -381 604 -369 608
rect -276 604 -264 608
rect -887 589 -875 593
rect -782 589 -770 593
rect -642 593 -630 597
rect -537 593 -525 597
rect -642 580 -630 584
rect -537 580 -525 584
rect -120 543 -116 555
rect -107 543 -103 555
rect -94 543 -90 555
rect -68 543 -64 555
rect -55 543 -51 555
rect -42 543 -38 555
rect 88 543 92 555
rect 101 543 105 555
rect 114 543 118 555
rect 140 543 144 555
rect 153 543 157 555
rect 166 543 170 555
rect -203 528 -199 540
rect -190 528 -186 540
rect -381 499 -369 503
rect -887 484 -875 488
rect -381 486 -369 490
rect -887 471 -875 475
rect -642 475 -630 479
rect -381 474 -369 478
rect -276 474 -264 478
rect -887 459 -875 463
rect -782 459 -770 463
rect -642 462 -630 466
rect -381 461 -369 465
rect -276 461 -264 465
rect -887 446 -875 450
rect -782 446 -770 450
rect -642 450 -630 454
rect -537 450 -525 454
rect -381 448 -369 452
rect -276 448 -264 452
rect -887 433 -875 437
rect -782 433 -770 437
rect -642 437 -630 441
rect -537 437 -525 441
rect -145 438 -141 450
rect -132 438 -128 450
rect -120 438 -116 450
rect -107 438 -103 450
rect -94 438 -90 450
rect -68 438 -64 450
rect -55 438 -51 450
rect -42 438 -38 450
rect 63 438 67 450
rect 76 438 80 450
rect 88 438 92 450
rect 101 438 105 450
rect 114 438 118 450
rect 140 438 144 450
rect 153 438 157 450
rect 166 438 170 450
rect -642 424 -630 428
rect -537 424 -525 428
rect -381 422 -369 426
rect -276 422 -264 426
rect -887 407 -875 411
rect -782 407 -770 411
rect -381 409 -369 413
rect -276 409 -264 413
rect -887 394 -875 398
rect -782 394 -770 398
rect -642 398 -630 402
rect -537 398 -525 402
rect -381 396 -369 400
rect -276 396 -264 400
rect -887 381 -875 385
rect -782 381 -770 385
rect -642 385 -630 389
rect -537 385 -525 389
rect -642 372 -630 376
rect -537 372 -525 376
rect 154 338 158 350
rect 167 338 171 350
rect 180 338 184 350
rect 206 338 210 350
rect 219 338 223 350
rect 232 338 236 350
rect 362 338 366 350
rect 375 338 379 350
rect 388 338 392 350
rect 414 338 418 350
rect 427 338 431 350
rect 440 338 444 350
rect 71 323 75 335
rect 84 323 88 335
rect -915 303 -903 307
rect -335 298 -331 318
rect -325 298 -321 318
rect -311 298 -307 318
rect -291 298 -287 318
rect -271 298 -267 318
rect -263 298 -259 318
rect -253 298 -249 318
rect -915 290 -903 294
rect -742 283 -738 295
rect -729 283 -725 295
rect -716 283 -712 295
rect -690 283 -686 295
rect -677 283 -673 295
rect -664 283 -660 295
rect -534 283 -530 295
rect -521 283 -517 295
rect -508 283 -504 295
rect -482 283 -478 295
rect -469 283 -465 295
rect -456 283 -452 295
rect -825 268 -821 280
rect -812 268 -808 280
rect -1005 245 -993 249
rect -1005 232 -993 236
rect -176 289 -172 296
rect -164 289 -160 296
rect -151 289 -147 296
rect -126 289 -122 296
rect -98 289 -94 296
rect -84 289 -80 296
rect -72 289 -68 296
rect -1005 220 -993 224
rect -900 220 -888 224
rect 129 233 133 245
rect 142 233 146 245
rect 154 233 158 245
rect 167 233 171 245
rect 180 233 184 245
rect 206 233 210 245
rect 219 233 223 245
rect 232 233 236 245
rect 337 233 341 245
rect 350 233 354 245
rect 362 233 366 245
rect 375 233 379 245
rect 388 233 392 245
rect 414 233 418 245
rect 427 233 431 245
rect 440 233 444 245
rect -1005 207 -993 211
rect -900 207 -888 211
rect -1005 194 -993 198
rect -900 194 -888 198
rect -335 190 -331 210
rect -325 190 -321 210
rect -315 190 -311 210
rect -307 190 -303 210
rect -297 190 -293 210
rect -767 178 -763 190
rect -754 178 -750 190
rect -742 178 -738 190
rect -729 178 -725 190
rect -716 178 -712 190
rect -690 178 -686 190
rect -677 178 -673 190
rect -664 178 -660 190
rect -559 178 -555 190
rect -546 178 -542 190
rect -534 178 -530 190
rect -521 178 -517 190
rect -508 178 -504 190
rect -482 178 -478 190
rect -469 178 -465 190
rect -456 178 -452 190
rect -1005 168 -993 172
rect -900 168 -888 172
rect -1005 155 -993 159
rect -900 155 -888 159
rect -1005 142 -993 146
rect -900 142 -888 146
rect -148 149 -143 160
rect -133 149 -129 160
rect -124 149 -120 160
rect -114 149 -110 160
rect -102 149 -98 160
rect -335 120 -331 140
rect -325 120 -321 140
rect -311 120 -307 140
rect -291 120 -287 140
rect -271 120 -267 140
rect -263 120 -259 140
rect -253 120 -249 140
rect -755 69 -751 81
rect -742 69 -738 81
rect -729 69 -725 81
rect -703 69 -699 81
rect -690 69 -686 81
rect -677 69 -673 81
rect -547 69 -543 81
rect -534 69 -530 81
rect -521 69 -517 81
rect -495 69 -491 81
rect -482 69 -478 81
rect -469 69 -465 81
rect -48 148 -42 159
rect -14 148 -9 159
rect -1 148 4 159
rect 12 148 16 159
rect 63 123 67 130
rect 75 123 79 130
rect 88 123 92 130
rect 113 123 117 130
rect 141 123 145 130
rect 155 123 159 130
rect 167 123 171 130
rect -838 54 -834 66
rect -825 54 -821 66
rect -1005 37 -993 41
rect -1005 24 -993 28
rect 375 111 379 123
rect 388 111 392 123
rect 401 111 405 123
rect 427 111 431 123
rect 440 111 444 123
rect 453 111 457 123
rect 583 111 587 123
rect 596 111 600 123
rect 609 111 613 123
rect 635 111 639 123
rect 648 111 652 123
rect 661 111 665 123
rect 292 96 296 108
rect 305 96 309 108
rect -1005 12 -993 16
rect -900 12 -888 16
rect -335 12 -331 32
rect -325 12 -321 32
rect -315 12 -311 32
rect -307 12 -303 32
rect -297 12 -293 32
rect -1005 -1 -993 3
rect -900 -1 -888 3
rect -173 7 -168 18
rect -158 7 -154 18
rect -149 7 -145 18
rect -139 7 -135 18
rect -127 7 -123 18
rect -1005 -14 -993 -10
rect -900 -14 -888 -10
rect -780 -36 -776 -24
rect -767 -36 -763 -24
rect -755 -36 -751 -24
rect -742 -36 -738 -24
rect -729 -36 -725 -24
rect -703 -36 -699 -24
rect -690 -36 -686 -24
rect -677 -36 -673 -24
rect -572 -36 -568 -24
rect -559 -36 -555 -24
rect -547 -36 -543 -24
rect -534 -36 -530 -24
rect -521 -36 -517 -24
rect -495 -36 -491 -24
rect -482 -36 -478 -24
rect -469 -36 -465 -24
rect 350 6 354 18
rect 363 6 367 18
rect 375 6 379 18
rect 388 6 392 18
rect 401 6 405 18
rect 427 6 431 18
rect 440 6 444 18
rect 453 6 457 18
rect 558 6 562 18
rect 571 6 575 18
rect 583 6 587 18
rect 596 6 600 18
rect 609 6 613 18
rect 635 6 639 18
rect 648 6 652 18
rect 661 6 665 18
rect -90 -7 -85 4
rect -75 -7 -71 4
rect -66 -7 -62 4
rect -56 -7 -52 4
rect -44 -7 -40 4
rect -1005 -40 -993 -36
rect -900 -40 -888 -36
rect -1005 -53 -993 -49
rect -900 -53 -888 -49
rect -1005 -66 -993 -62
rect -900 -66 -888 -62
rect -335 -58 -331 -38
rect -325 -58 -321 -38
rect -311 -58 -307 -38
rect -291 -58 -287 -38
rect -271 -58 -267 -38
rect -263 -58 -259 -38
rect -253 -58 -249 -38
rect 11 -39 17 -28
rect 45 -39 50 -28
rect 58 -39 63 -28
rect 71 -39 75 -28
rect 123 -38 127 -31
rect 135 -38 139 -31
rect 148 -38 152 -31
rect 173 -38 177 -31
rect 201 -38 205 -31
rect 215 -38 219 -31
rect 227 -38 231 -31
rect -182 -91 -177 -80
rect -167 -91 -163 -80
rect -158 -91 -154 -80
rect -148 -91 -144 -80
rect -136 -91 -132 -80
rect -90 -112 -84 -101
rect -56 -112 -51 -101
rect -43 -112 -38 -101
rect -30 -112 -26 -101
rect 369 -103 373 -91
rect 382 -103 386 -91
rect 395 -103 399 -91
rect 421 -103 425 -91
rect 434 -103 438 -91
rect 447 -103 451 -91
rect 577 -103 581 -91
rect 590 -103 594 -91
rect 603 -103 607 -91
rect 629 -103 633 -91
rect 642 -103 646 -91
rect 655 -103 659 -91
rect -757 -162 -753 -150
rect -744 -162 -740 -150
rect -731 -162 -727 -150
rect -705 -162 -701 -150
rect -692 -162 -688 -150
rect -679 -162 -675 -150
rect -549 -162 -545 -150
rect -536 -162 -532 -150
rect -523 -162 -519 -150
rect -497 -162 -493 -150
rect -484 -162 -480 -150
rect -471 -162 -467 -150
rect -840 -177 -836 -165
rect -827 -177 -823 -165
rect -335 -166 -331 -146
rect -325 -166 -321 -146
rect -315 -166 -311 -146
rect -307 -166 -303 -146
rect -297 -166 -293 -146
rect 286 -118 290 -106
rect 299 -118 303 -106
rect -154 -210 -149 -199
rect -139 -210 -135 -199
rect -130 -210 -126 -199
rect -120 -210 -116 -199
rect -108 -210 -104 -199
rect 344 -208 348 -196
rect 357 -208 361 -196
rect 369 -208 373 -196
rect 382 -208 386 -196
rect 395 -208 399 -196
rect 421 -208 425 -196
rect 434 -208 438 -196
rect 447 -208 451 -196
rect 552 -208 556 -196
rect 565 -208 569 -196
rect 577 -208 581 -196
rect 590 -208 594 -196
rect 603 -208 607 -196
rect 629 -208 633 -196
rect 642 -208 646 -196
rect 655 -208 659 -196
rect -335 -236 -331 -216
rect -325 -236 -321 -216
rect -311 -236 -307 -216
rect -291 -236 -287 -216
rect -271 -236 -267 -216
rect -263 -236 -259 -216
rect -253 -236 -249 -216
rect -782 -267 -778 -255
rect -769 -267 -765 -255
rect -757 -267 -753 -255
rect -744 -267 -740 -255
rect -731 -267 -727 -255
rect -705 -267 -701 -255
rect -692 -267 -688 -255
rect -679 -267 -675 -255
rect -574 -267 -570 -255
rect -561 -267 -557 -255
rect -549 -267 -545 -255
rect -536 -267 -532 -255
rect -523 -267 -519 -255
rect -497 -267 -493 -255
rect -484 -267 -480 -255
rect -471 -267 -467 -255
rect -71 -224 -66 -213
rect -56 -224 -52 -213
rect -47 -224 -43 -213
rect -37 -224 -33 -213
rect -25 -224 -21 -213
rect 12 -232 17 -221
rect 27 -232 31 -221
rect 36 -232 40 -221
rect 46 -232 50 -221
rect 58 -232 62 -221
rect 91 -275 97 -264
rect 125 -275 130 -264
rect 138 -275 143 -264
rect 151 -275 155 -264
rect -335 -344 -331 -324
rect -325 -344 -321 -324
rect -315 -344 -311 -324
rect -307 -344 -303 -324
rect -297 -344 -293 -324
rect -139 -326 -134 -315
rect -124 -326 -120 -315
rect -115 -326 -111 -315
rect -105 -326 -101 -315
rect -93 -326 -89 -315
rect -766 -377 -762 -365
rect -753 -377 -749 -365
rect -740 -377 -736 -365
rect -714 -377 -710 -365
rect -701 -377 -697 -365
rect -688 -377 -684 -365
rect -558 -377 -554 -365
rect -545 -377 -541 -365
rect -532 -377 -528 -365
rect -506 -377 -502 -365
rect -493 -377 -489 -365
rect -480 -377 -476 -365
rect 282 -327 286 -315
rect 295 -327 299 -315
rect 308 -327 312 -315
rect 334 -327 338 -315
rect 347 -327 351 -315
rect 360 -327 364 -315
rect 490 -327 494 -315
rect 503 -327 507 -315
rect 516 -327 520 -315
rect 542 -327 546 -315
rect 555 -327 559 -315
rect 568 -327 572 -315
rect -56 -340 -51 -329
rect -41 -340 -37 -329
rect -32 -340 -28 -329
rect -22 -340 -18 -329
rect -10 -340 -6 -329
rect -849 -392 -845 -380
rect -836 -392 -832 -380
rect 199 -342 203 -330
rect 212 -342 216 -330
rect 55 -392 61 -381
rect 89 -392 94 -381
rect 102 -392 107 -381
rect 115 -392 119 -381
rect -141 -420 -136 -409
rect -126 -420 -122 -409
rect -117 -420 -113 -409
rect -107 -420 -103 -409
rect -95 -420 -91 -409
rect -46 -435 -40 -424
rect -12 -435 -7 -424
rect 1 -435 6 -424
rect 14 -435 18 -424
rect -791 -482 -787 -470
rect -778 -482 -774 -470
rect -766 -482 -762 -470
rect -753 -482 -749 -470
rect -740 -482 -736 -470
rect -714 -482 -710 -470
rect -701 -482 -697 -470
rect -688 -482 -684 -470
rect -583 -482 -579 -470
rect -570 -482 -566 -470
rect -558 -482 -554 -470
rect -545 -482 -541 -470
rect -532 -482 -528 -470
rect -506 -482 -502 -470
rect -493 -482 -489 -470
rect -480 -482 -476 -470
rect 257 -432 261 -420
rect 270 -432 274 -420
rect 282 -432 286 -420
rect 295 -432 299 -420
rect 308 -432 312 -420
rect 334 -432 338 -420
rect 347 -432 351 -420
rect 360 -432 364 -420
rect 465 -432 469 -420
rect 478 -432 482 -420
rect 490 -432 494 -420
rect 503 -432 507 -420
rect 516 -432 520 -420
rect 542 -432 546 -420
rect 555 -432 559 -420
rect 568 -432 572 -420
<< polysilicon >>
rect -328 760 -325 762
rect -318 760 -291 762
rect -279 760 -276 762
rect -834 745 -831 747
rect -824 745 -797 747
rect -785 745 -782 747
rect -589 736 -586 738
rect -579 736 -552 738
rect -540 736 -537 738
rect -418 702 -415 704
rect -408 702 -381 704
rect -369 702 -366 704
rect -924 687 -921 689
rect -914 687 -887 689
rect -875 687 -872 689
rect -679 678 -676 680
rect -669 678 -642 680
rect -630 678 -627 680
rect -443 677 -440 679
rect -434 677 -381 679
rect -369 677 -366 679
rect -338 677 -335 679
rect -329 677 -276 679
rect -264 677 -261 679
rect -949 662 -946 664
rect -940 662 -887 664
rect -875 662 -872 664
rect -844 662 -841 664
rect -835 662 -782 664
rect -770 662 -767 664
rect -443 662 -440 664
rect -434 662 -381 664
rect -369 662 -366 664
rect -338 662 -335 664
rect -329 662 -276 664
rect -264 662 -261 664
rect -704 653 -701 655
rect -695 653 -642 655
rect -630 653 -627 655
rect -599 653 -596 655
rect -590 653 -537 655
rect -525 653 -522 655
rect -949 647 -946 649
rect -940 647 -887 649
rect -875 647 -872 649
rect -844 647 -841 649
rect -835 647 -782 649
rect -770 647 -767 649
rect -704 638 -701 640
rect -695 638 -642 640
rect -630 638 -627 640
rect -599 638 -596 640
rect -590 638 -537 640
rect -525 638 -522 640
rect -443 625 -440 627
rect -434 625 -381 627
rect -369 625 -366 627
rect -338 625 -335 627
rect -329 625 -276 627
rect -264 625 -261 627
rect -949 610 -946 612
rect -940 610 -887 612
rect -875 610 -872 612
rect -844 610 -841 612
rect -835 610 -782 612
rect -770 610 -767 612
rect -443 610 -440 612
rect -434 610 -381 612
rect -369 610 -366 612
rect -338 610 -335 612
rect -329 610 -276 612
rect -264 610 -261 612
rect -704 601 -701 603
rect -695 601 -642 603
rect -630 601 -627 603
rect -599 601 -596 603
rect -590 601 -537 603
rect -525 601 -522 603
rect -949 595 -946 597
rect -940 595 -887 597
rect -875 595 -872 597
rect -844 595 -841 597
rect -835 595 -782 597
rect -770 595 -767 597
rect -704 586 -701 588
rect -695 586 -642 588
rect -630 586 -627 588
rect -599 586 -596 588
rect -590 586 -537 588
rect -525 586 -522 588
rect -113 555 -111 558
rect -98 555 -96 558
rect -61 555 -59 558
rect -46 555 -44 558
rect 95 555 97 558
rect 110 555 112 558
rect 147 555 149 558
rect 162 555 164 558
rect -196 540 -194 543
rect -196 501 -194 528
rect -418 494 -415 496
rect -408 494 -381 496
rect -369 494 -366 496
rect -196 491 -194 494
rect -113 490 -111 543
rect -98 490 -96 543
rect -61 490 -59 543
rect -46 490 -44 543
rect 95 490 97 543
rect 110 490 112 543
rect 147 490 149 543
rect 162 490 164 543
rect -113 481 -111 484
rect -98 481 -96 484
rect -61 481 -59 484
rect -46 481 -44 484
rect 95 481 97 484
rect 110 481 112 484
rect 147 481 149 484
rect 162 481 164 484
rect -924 479 -921 481
rect -914 479 -887 481
rect -875 479 -872 481
rect -679 470 -676 472
rect -669 470 -642 472
rect -630 470 -627 472
rect -443 469 -440 471
rect -434 469 -381 471
rect -369 469 -366 471
rect -338 469 -335 471
rect -329 469 -276 471
rect -264 469 -261 471
rect -949 454 -946 456
rect -940 454 -887 456
rect -875 454 -872 456
rect -844 454 -841 456
rect -835 454 -782 456
rect -770 454 -767 456
rect -443 454 -440 456
rect -434 454 -381 456
rect -369 454 -366 456
rect -338 454 -335 456
rect -329 454 -276 456
rect -264 454 -261 456
rect -138 450 -136 453
rect -113 450 -111 453
rect -98 450 -96 453
rect -61 450 -59 453
rect -46 450 -44 453
rect 70 450 72 453
rect 95 450 97 453
rect 110 450 112 453
rect 147 450 149 453
rect 162 450 164 453
rect -704 445 -701 447
rect -695 445 -642 447
rect -630 445 -627 447
rect -599 445 -596 447
rect -590 445 -537 447
rect -525 445 -522 447
rect -949 439 -946 441
rect -940 439 -887 441
rect -875 439 -872 441
rect -844 439 -841 441
rect -835 439 -782 441
rect -770 439 -767 441
rect -704 430 -701 432
rect -695 430 -642 432
rect -630 430 -627 432
rect -599 430 -596 432
rect -590 430 -537 432
rect -525 430 -522 432
rect -443 417 -440 419
rect -434 417 -381 419
rect -369 417 -366 419
rect -338 417 -335 419
rect -329 417 -276 419
rect -264 417 -261 419
rect -138 411 -136 438
rect -949 402 -946 404
rect -940 402 -887 404
rect -875 402 -872 404
rect -844 402 -841 404
rect -835 402 -782 404
rect -770 402 -767 404
rect -443 402 -440 404
rect -434 402 -381 404
rect -369 402 -366 404
rect -338 402 -335 404
rect -329 402 -276 404
rect -264 402 -261 404
rect -138 401 -136 404
rect -704 393 -701 395
rect -695 393 -642 395
rect -630 393 -627 395
rect -599 393 -596 395
rect -590 393 -537 395
rect -525 393 -522 395
rect -949 387 -946 389
rect -940 387 -887 389
rect -875 387 -872 389
rect -844 387 -841 389
rect -835 387 -782 389
rect -770 387 -767 389
rect -113 385 -111 438
rect -98 385 -96 438
rect -61 385 -59 438
rect -46 385 -44 438
rect 70 411 72 438
rect 70 401 72 404
rect 95 385 97 438
rect 110 385 112 438
rect 147 385 149 438
rect 162 385 164 438
rect -704 378 -701 380
rect -695 378 -642 380
rect -630 378 -627 380
rect -599 378 -596 380
rect -590 378 -537 380
rect -525 378 -522 380
rect -113 376 -111 379
rect -98 376 -96 379
rect -61 376 -59 379
rect -46 376 -44 379
rect 95 376 97 379
rect 110 376 112 379
rect 147 376 149 379
rect 162 376 164 379
rect 161 350 163 353
rect 176 350 178 353
rect 213 350 215 353
rect 228 350 230 353
rect 369 350 371 353
rect 384 350 386 353
rect 421 350 423 353
rect 436 350 438 353
rect 78 335 80 338
rect -329 318 -327 321
rect -305 318 -303 321
rect -295 318 -293 321
rect -285 318 -283 321
rect -275 318 -273 321
rect -257 318 -255 321
rect -952 298 -949 300
rect -942 298 -915 300
rect -903 298 -900 300
rect -735 295 -733 298
rect -720 295 -718 298
rect -683 295 -681 298
rect -668 295 -666 298
rect -527 295 -525 298
rect -512 295 -510 298
rect -475 295 -473 298
rect -460 295 -458 298
rect -329 285 -327 298
rect -818 280 -816 283
rect -1042 240 -1039 242
rect -1032 240 -1005 242
rect -993 240 -990 242
rect -818 241 -816 268
rect -818 231 -816 234
rect -735 230 -733 283
rect -720 230 -718 283
rect -683 230 -681 283
rect -668 230 -666 283
rect -527 230 -525 283
rect -512 230 -510 283
rect -475 230 -473 283
rect -460 230 -458 283
rect -329 272 -327 275
rect -305 250 -303 298
rect -295 250 -293 298
rect -285 250 -283 298
rect -275 250 -273 298
rect -257 285 -255 298
rect -169 296 -167 299
rect -144 296 -142 299
rect -132 296 -130 299
rect -118 296 -116 299
rect -105 296 -103 299
rect -77 296 -75 299
rect 78 296 80 323
rect -257 272 -255 275
rect -169 259 -167 289
rect -169 247 -167 250
rect -305 237 -303 240
rect -295 237 -293 240
rect -285 237 -283 240
rect -275 237 -273 240
rect -735 221 -733 224
rect -720 221 -718 224
rect -683 221 -681 224
rect -668 221 -666 224
rect -527 221 -525 224
rect -512 221 -510 224
rect -475 221 -473 224
rect -460 221 -458 224
rect -144 223 -142 289
rect -132 223 -130 289
rect -118 223 -116 289
rect -105 223 -103 289
rect -77 260 -75 289
rect 78 286 80 289
rect 161 285 163 338
rect 176 285 178 338
rect 213 285 215 338
rect 228 285 230 338
rect 369 285 371 338
rect 384 285 386 338
rect 421 285 423 338
rect 436 285 438 338
rect 161 276 163 279
rect 176 276 178 279
rect 213 276 215 279
rect 228 276 230 279
rect 369 276 371 279
rect 384 276 386 279
rect 421 276 423 279
rect 436 276 438 279
rect -77 247 -75 251
rect 136 245 138 248
rect 161 245 163 248
rect 176 245 178 248
rect 213 245 215 248
rect 228 245 230 248
rect 344 245 346 248
rect 369 245 371 248
rect 384 245 386 248
rect 421 245 423 248
rect 436 245 438 248
rect -1067 215 -1064 217
rect -1058 215 -1005 217
rect -993 215 -990 217
rect -962 215 -959 217
rect -953 215 -900 217
rect -888 215 -885 217
rect -329 210 -327 213
rect -319 210 -317 213
rect -301 210 -299 213
rect -144 210 -142 213
rect -132 210 -130 213
rect -118 210 -116 213
rect -105 210 -103 213
rect -1067 200 -1064 202
rect -1058 200 -1005 202
rect -993 200 -990 202
rect -962 200 -959 202
rect -953 200 -900 202
rect -888 200 -885 202
rect -760 190 -758 193
rect -735 190 -733 193
rect -720 190 -718 193
rect -683 190 -681 193
rect -668 190 -666 193
rect -552 190 -550 193
rect -527 190 -525 193
rect -512 190 -510 193
rect -475 190 -473 193
rect -460 190 -458 193
rect 136 206 138 233
rect 136 196 138 199
rect -1067 163 -1064 165
rect -1058 163 -1005 165
rect -993 163 -990 165
rect -962 163 -959 165
rect -953 163 -900 165
rect -888 163 -885 165
rect -760 151 -758 178
rect -1067 148 -1064 150
rect -1058 148 -1005 150
rect -993 148 -990 150
rect -962 148 -959 150
rect -953 148 -900 150
rect -888 148 -885 150
rect -760 141 -758 144
rect -735 125 -733 178
rect -720 125 -718 178
rect -683 125 -681 178
rect -668 125 -666 178
rect -552 151 -550 178
rect -552 141 -550 144
rect -527 125 -525 178
rect -512 125 -510 178
rect -475 125 -473 178
rect -460 125 -458 178
rect -329 170 -327 190
rect -319 170 -317 190
rect -301 170 -299 190
rect 161 180 163 233
rect 176 180 178 233
rect 213 180 215 233
rect 228 180 230 233
rect 344 206 346 233
rect 344 196 346 199
rect 369 180 371 233
rect 384 180 386 233
rect 421 180 423 233
rect 436 180 438 233
rect 161 171 163 174
rect 176 171 178 174
rect 213 171 215 174
rect 228 171 230 174
rect 369 171 371 174
rect 384 171 386 174
rect 421 171 423 174
rect 436 171 438 174
rect -141 160 -139 163
rect -128 160 -126 163
rect -106 160 -104 163
rect -329 157 -327 160
rect -319 157 -317 160
rect -301 157 -299 160
rect -38 159 -36 163
rect -20 159 -18 163
rect 7 159 9 162
rect -329 140 -327 143
rect -305 140 -303 143
rect -295 140 -293 143
rect -285 140 -283 143
rect -275 140 -273 143
rect -257 140 -255 143
rect -735 116 -733 119
rect -720 116 -718 119
rect -683 116 -681 119
rect -668 116 -666 119
rect -527 116 -525 119
rect -512 116 -510 119
rect -475 116 -473 119
rect -460 116 -458 119
rect -329 107 -327 120
rect -329 94 -327 97
rect -748 81 -746 84
rect -733 81 -731 84
rect -696 81 -694 84
rect -681 81 -679 84
rect -540 81 -538 84
rect -525 81 -523 84
rect -488 81 -486 84
rect -473 81 -471 84
rect -305 72 -303 120
rect -295 72 -293 120
rect -285 72 -283 120
rect -275 72 -273 120
rect -257 107 -255 120
rect -141 108 -139 149
rect -128 108 -126 149
rect -106 109 -104 149
rect -141 97 -139 100
rect -128 97 -126 100
rect -106 98 -104 101
rect -257 94 -255 97
rect -38 95 -36 148
rect -20 95 -18 148
rect 7 95 9 148
rect 70 130 72 133
rect 95 130 97 133
rect 107 130 109 133
rect 121 130 123 133
rect 134 130 136 133
rect 162 130 164 133
rect 382 123 384 126
rect 397 123 399 126
rect 434 123 436 126
rect 449 123 451 126
rect 590 123 592 126
rect 605 123 607 126
rect 642 123 644 126
rect 657 123 659 126
rect 70 93 72 123
rect -38 84 -36 87
rect -20 84 -18 87
rect 7 84 9 87
rect 70 81 72 84
rect -831 66 -829 69
rect -1042 32 -1039 34
rect -1032 32 -1005 34
rect -993 32 -990 34
rect -831 27 -829 54
rect -831 17 -829 20
rect -748 16 -746 69
rect -733 16 -731 69
rect -696 16 -694 69
rect -681 16 -679 69
rect -540 16 -538 69
rect -525 16 -523 69
rect -488 16 -486 69
rect -473 16 -471 69
rect -305 59 -303 62
rect -295 59 -293 62
rect -285 59 -283 62
rect -275 59 -273 62
rect 95 57 97 123
rect 107 57 109 123
rect 121 57 123 123
rect 134 57 136 123
rect 162 94 164 123
rect 299 108 301 111
rect 162 81 164 85
rect 299 69 301 96
rect 299 59 301 62
rect 382 58 384 111
rect 397 58 399 111
rect 434 58 436 111
rect 449 58 451 111
rect 590 58 592 111
rect 605 58 607 111
rect 642 58 644 111
rect 657 58 659 111
rect 382 49 384 52
rect 397 49 399 52
rect 434 49 436 52
rect 449 49 451 52
rect 590 49 592 52
rect 605 49 607 52
rect 642 49 644 52
rect 657 49 659 52
rect 95 44 97 47
rect 107 44 109 47
rect 121 44 123 47
rect 134 44 136 47
rect -329 32 -327 35
rect -319 32 -317 35
rect -301 32 -299 35
rect -166 18 -164 21
rect -153 18 -151 21
rect -131 18 -129 21
rect 357 18 359 21
rect 382 18 384 21
rect 397 18 399 21
rect 434 18 436 21
rect 449 18 451 21
rect 565 18 567 21
rect 590 18 592 21
rect 605 18 607 21
rect 642 18 644 21
rect 657 18 659 21
rect -1067 7 -1064 9
rect -1058 7 -1005 9
rect -993 7 -990 9
rect -962 7 -959 9
rect -953 7 -900 9
rect -888 7 -885 9
rect -748 7 -746 10
rect -733 7 -731 10
rect -696 7 -694 10
rect -681 7 -679 10
rect -540 7 -538 10
rect -525 7 -523 10
rect -488 7 -486 10
rect -473 7 -471 10
rect -1067 -8 -1064 -6
rect -1058 -8 -1005 -6
rect -993 -8 -990 -6
rect -962 -8 -959 -6
rect -953 -8 -900 -6
rect -888 -8 -885 -6
rect -329 -8 -327 12
rect -319 -8 -317 12
rect -301 -8 -299 12
rect -329 -21 -327 -18
rect -319 -21 -317 -18
rect -301 -21 -299 -18
rect -773 -24 -771 -21
rect -748 -24 -746 -21
rect -733 -24 -731 -21
rect -696 -24 -694 -21
rect -681 -24 -679 -21
rect -565 -24 -563 -21
rect -540 -24 -538 -21
rect -525 -24 -523 -21
rect -488 -24 -486 -21
rect -473 -24 -471 -21
rect -166 -34 -164 7
rect -153 -34 -151 7
rect -131 -33 -129 7
rect -83 4 -81 7
rect -70 4 -68 7
rect -48 4 -46 7
rect -1067 -45 -1064 -43
rect -1058 -45 -1005 -43
rect -993 -45 -990 -43
rect -962 -45 -959 -43
rect -953 -45 -900 -43
rect -888 -45 -885 -43
rect -1067 -60 -1064 -58
rect -1058 -60 -1005 -58
rect -993 -60 -990 -58
rect -962 -60 -959 -58
rect -953 -60 -900 -58
rect -888 -60 -885 -58
rect -773 -63 -771 -36
rect -773 -73 -771 -70
rect -748 -89 -746 -36
rect -733 -89 -731 -36
rect -696 -89 -694 -36
rect -681 -89 -679 -36
rect -565 -63 -563 -36
rect -565 -73 -563 -70
rect -540 -89 -538 -36
rect -525 -89 -523 -36
rect -488 -89 -486 -36
rect -473 -89 -471 -36
rect -329 -38 -327 -35
rect -305 -38 -303 -35
rect -295 -38 -293 -35
rect -285 -38 -283 -35
rect -275 -38 -273 -35
rect -257 -38 -255 -35
rect -166 -45 -164 -42
rect -153 -45 -151 -42
rect -131 -44 -129 -41
rect -83 -48 -81 -7
rect -70 -48 -68 -7
rect -48 -47 -46 -7
rect 357 -21 359 6
rect 21 -28 23 -24
rect 39 -28 41 -24
rect 66 -28 68 -25
rect 130 -31 132 -28
rect 155 -31 157 -28
rect 167 -31 169 -28
rect 181 -31 183 -28
rect 194 -31 196 -28
rect 222 -31 224 -28
rect 357 -31 359 -28
rect -329 -71 -327 -58
rect -329 -84 -327 -81
rect -748 -98 -746 -95
rect -733 -98 -731 -95
rect -696 -98 -694 -95
rect -681 -98 -679 -95
rect -540 -98 -538 -95
rect -525 -98 -523 -95
rect -488 -98 -486 -95
rect -473 -98 -471 -95
rect -305 -106 -303 -58
rect -295 -106 -293 -58
rect -285 -106 -283 -58
rect -275 -106 -273 -58
rect -257 -71 -255 -58
rect -83 -59 -81 -56
rect -70 -59 -68 -56
rect -48 -58 -46 -55
rect -175 -80 -173 -77
rect -162 -80 -160 -77
rect -140 -80 -138 -77
rect -257 -84 -255 -81
rect -305 -119 -303 -116
rect -295 -119 -293 -116
rect -285 -119 -283 -116
rect -275 -119 -273 -116
rect -175 -132 -173 -91
rect -162 -132 -160 -91
rect -140 -131 -138 -91
rect 21 -92 23 -39
rect 39 -92 41 -39
rect 66 -92 68 -39
rect 130 -68 132 -38
rect 130 -80 132 -77
rect -80 -101 -78 -97
rect -62 -101 -60 -97
rect -35 -101 -33 -98
rect 21 -103 23 -100
rect 39 -103 41 -100
rect 66 -103 68 -100
rect 155 -104 157 -38
rect 167 -104 169 -38
rect 181 -104 183 -38
rect 194 -104 196 -38
rect 222 -67 224 -38
rect 382 -47 384 6
rect 397 -47 399 6
rect 434 -47 436 6
rect 449 -47 451 6
rect 565 -21 567 6
rect 565 -31 567 -28
rect 590 -47 592 6
rect 605 -47 607 6
rect 642 -47 644 6
rect 657 -47 659 6
rect 382 -56 384 -53
rect 397 -56 399 -53
rect 434 -56 436 -53
rect 449 -56 451 -53
rect 590 -56 592 -53
rect 605 -56 607 -53
rect 642 -56 644 -53
rect 657 -56 659 -53
rect 222 -80 224 -76
rect 376 -91 378 -88
rect 391 -91 393 -88
rect 428 -91 430 -88
rect 443 -91 445 -88
rect 584 -91 586 -88
rect 599 -91 601 -88
rect 636 -91 638 -88
rect 651 -91 653 -88
rect -175 -143 -173 -140
rect -162 -143 -160 -140
rect -140 -142 -138 -139
rect -329 -146 -327 -143
rect -319 -146 -317 -143
rect -301 -146 -299 -143
rect -750 -150 -748 -147
rect -735 -150 -733 -147
rect -698 -150 -696 -147
rect -683 -150 -681 -147
rect -542 -150 -540 -147
rect -527 -150 -525 -147
rect -490 -150 -488 -147
rect -475 -150 -473 -147
rect -833 -165 -831 -162
rect -833 -204 -831 -177
rect -833 -214 -831 -211
rect -750 -215 -748 -162
rect -735 -215 -733 -162
rect -698 -215 -696 -162
rect -683 -215 -681 -162
rect -542 -215 -540 -162
rect -527 -215 -525 -162
rect -490 -215 -488 -162
rect -475 -215 -473 -162
rect -80 -165 -78 -112
rect -62 -165 -60 -112
rect -35 -165 -33 -112
rect 293 -106 295 -103
rect 155 -117 157 -114
rect 167 -117 169 -114
rect 181 -117 183 -114
rect 194 -117 196 -114
rect 293 -145 295 -118
rect 293 -155 295 -152
rect 376 -156 378 -103
rect 391 -156 393 -103
rect 428 -156 430 -103
rect 443 -156 445 -103
rect 584 -156 586 -103
rect 599 -156 601 -103
rect 636 -156 638 -103
rect 651 -156 653 -103
rect 376 -165 378 -162
rect 391 -165 393 -162
rect 428 -165 430 -162
rect 443 -165 445 -162
rect 584 -165 586 -162
rect 599 -165 601 -162
rect 636 -165 638 -162
rect 651 -165 653 -162
rect -329 -186 -327 -166
rect -319 -186 -317 -166
rect -301 -186 -299 -166
rect -80 -176 -78 -173
rect -62 -176 -60 -173
rect -35 -176 -33 -173
rect 351 -196 353 -193
rect 376 -196 378 -193
rect 391 -196 393 -193
rect 428 -196 430 -193
rect 443 -196 445 -193
rect 559 -196 561 -193
rect 584 -196 586 -193
rect 599 -196 601 -193
rect 636 -196 638 -193
rect 651 -196 653 -193
rect -329 -199 -327 -196
rect -319 -199 -317 -196
rect -301 -199 -299 -196
rect -147 -199 -145 -196
rect -134 -199 -132 -196
rect -112 -199 -110 -196
rect -329 -216 -327 -213
rect -305 -216 -303 -213
rect -295 -216 -293 -213
rect -285 -216 -283 -213
rect -275 -216 -273 -213
rect -257 -216 -255 -213
rect -750 -224 -748 -221
rect -735 -224 -733 -221
rect -698 -224 -696 -221
rect -683 -224 -681 -221
rect -542 -224 -540 -221
rect -527 -224 -525 -221
rect -490 -224 -488 -221
rect -475 -224 -473 -221
rect -329 -249 -327 -236
rect -775 -255 -773 -252
rect -750 -255 -748 -252
rect -735 -255 -733 -252
rect -698 -255 -696 -252
rect -683 -255 -681 -252
rect -567 -255 -565 -252
rect -542 -255 -540 -252
rect -527 -255 -525 -252
rect -490 -255 -488 -252
rect -475 -255 -473 -252
rect -329 -262 -327 -259
rect -775 -294 -773 -267
rect -775 -304 -773 -301
rect -750 -320 -748 -267
rect -735 -320 -733 -267
rect -698 -320 -696 -267
rect -683 -320 -681 -267
rect -567 -294 -565 -267
rect -567 -304 -565 -301
rect -542 -320 -540 -267
rect -527 -320 -525 -267
rect -490 -320 -488 -267
rect -475 -320 -473 -267
rect -305 -284 -303 -236
rect -295 -284 -293 -236
rect -285 -284 -283 -236
rect -275 -284 -273 -236
rect -257 -249 -255 -236
rect -147 -251 -145 -210
rect -134 -251 -132 -210
rect -112 -250 -110 -210
rect -64 -213 -62 -210
rect -51 -213 -49 -210
rect -29 -213 -27 -210
rect 19 -221 21 -218
rect 32 -221 34 -218
rect 54 -221 56 -218
rect -257 -262 -255 -259
rect -147 -262 -145 -259
rect -134 -262 -132 -259
rect -112 -261 -110 -258
rect -64 -265 -62 -224
rect -51 -265 -49 -224
rect -29 -264 -27 -224
rect -64 -276 -62 -273
rect -51 -276 -49 -273
rect -29 -275 -27 -272
rect 19 -273 21 -232
rect 32 -273 34 -232
rect 54 -272 56 -232
rect 351 -235 353 -208
rect 351 -245 353 -242
rect 101 -264 103 -260
rect 119 -264 121 -260
rect 376 -261 378 -208
rect 391 -261 393 -208
rect 428 -261 430 -208
rect 443 -261 445 -208
rect 559 -235 561 -208
rect 559 -245 561 -242
rect 584 -261 586 -208
rect 599 -261 601 -208
rect 636 -261 638 -208
rect 651 -261 653 -208
rect 146 -264 148 -261
rect 376 -270 378 -267
rect 391 -270 393 -267
rect 428 -270 430 -267
rect 443 -270 445 -267
rect 584 -270 586 -267
rect 599 -270 601 -267
rect 636 -270 638 -267
rect 651 -270 653 -267
rect 19 -284 21 -281
rect 32 -284 34 -281
rect 54 -283 56 -280
rect -305 -297 -303 -294
rect -295 -297 -293 -294
rect -285 -297 -283 -294
rect -275 -297 -273 -294
rect -132 -315 -130 -312
rect -119 -315 -117 -312
rect -97 -315 -95 -312
rect -329 -324 -327 -321
rect -319 -324 -317 -321
rect -301 -324 -299 -321
rect -750 -329 -748 -326
rect -735 -329 -733 -326
rect -698 -329 -696 -326
rect -683 -329 -681 -326
rect -542 -329 -540 -326
rect -527 -329 -525 -326
rect -490 -329 -488 -326
rect -475 -329 -473 -326
rect -759 -365 -757 -362
rect -744 -365 -742 -362
rect -707 -365 -705 -362
rect -692 -365 -690 -362
rect -551 -365 -549 -362
rect -536 -365 -534 -362
rect -499 -365 -497 -362
rect -484 -365 -482 -362
rect -329 -364 -327 -344
rect -319 -364 -317 -344
rect -301 -364 -299 -344
rect -132 -367 -130 -326
rect -119 -367 -117 -326
rect -97 -366 -95 -326
rect -49 -329 -47 -326
rect -36 -329 -34 -326
rect -14 -329 -12 -326
rect 101 -328 103 -275
rect 119 -328 121 -275
rect 146 -328 148 -275
rect 289 -315 291 -312
rect 304 -315 306 -312
rect 341 -315 343 -312
rect 356 -315 358 -312
rect 497 -315 499 -312
rect 512 -315 514 -312
rect 549 -315 551 -312
rect 564 -315 566 -312
rect 206 -330 208 -327
rect 101 -339 103 -336
rect 119 -339 121 -336
rect 146 -339 148 -336
rect -329 -377 -327 -374
rect -319 -377 -317 -374
rect -301 -377 -299 -374
rect -842 -380 -840 -377
rect -842 -419 -840 -392
rect -842 -429 -840 -426
rect -759 -430 -757 -377
rect -744 -430 -742 -377
rect -707 -430 -705 -377
rect -692 -430 -690 -377
rect -551 -430 -549 -377
rect -536 -430 -534 -377
rect -499 -430 -497 -377
rect -484 -430 -482 -377
rect -132 -378 -130 -375
rect -119 -378 -117 -375
rect -97 -377 -95 -374
rect -49 -381 -47 -340
rect -36 -381 -34 -340
rect -14 -380 -12 -340
rect 206 -369 208 -342
rect 65 -381 67 -377
rect 83 -381 85 -377
rect 110 -381 112 -378
rect 206 -379 208 -376
rect 289 -380 291 -327
rect 304 -380 306 -327
rect 341 -380 343 -327
rect 356 -380 358 -327
rect 497 -380 499 -327
rect 512 -380 514 -327
rect 549 -380 551 -327
rect 564 -380 566 -327
rect -49 -392 -47 -389
rect -36 -392 -34 -389
rect -14 -391 -12 -388
rect 289 -389 291 -386
rect 304 -389 306 -386
rect 341 -389 343 -386
rect 356 -389 358 -386
rect 497 -389 499 -386
rect 512 -389 514 -386
rect 549 -389 551 -386
rect 564 -389 566 -386
rect -134 -409 -132 -406
rect -121 -409 -119 -406
rect -99 -409 -97 -406
rect -759 -439 -757 -436
rect -744 -439 -742 -436
rect -707 -439 -705 -436
rect -692 -439 -690 -436
rect -551 -439 -549 -436
rect -536 -439 -534 -436
rect -499 -439 -497 -436
rect -484 -439 -482 -436
rect -134 -461 -132 -420
rect -121 -461 -119 -420
rect -99 -460 -97 -420
rect -36 -424 -34 -420
rect -18 -424 -16 -420
rect 9 -424 11 -421
rect -784 -470 -782 -467
rect -759 -470 -757 -467
rect -744 -470 -742 -467
rect -707 -470 -705 -467
rect -692 -470 -690 -467
rect -576 -470 -574 -467
rect -551 -470 -549 -467
rect -536 -470 -534 -467
rect -499 -470 -497 -467
rect -484 -470 -482 -467
rect -134 -472 -132 -469
rect -121 -472 -119 -469
rect -99 -471 -97 -468
rect -784 -509 -782 -482
rect -784 -519 -782 -516
rect -759 -535 -757 -482
rect -744 -535 -742 -482
rect -707 -535 -705 -482
rect -692 -535 -690 -482
rect -576 -509 -574 -482
rect -576 -519 -574 -516
rect -551 -535 -549 -482
rect -536 -535 -534 -482
rect -499 -535 -497 -482
rect -484 -535 -482 -482
rect -36 -488 -34 -435
rect -18 -488 -16 -435
rect 9 -488 11 -435
rect 65 -445 67 -392
rect 83 -445 85 -392
rect 110 -445 112 -392
rect 264 -420 266 -417
rect 289 -420 291 -417
rect 304 -420 306 -417
rect 341 -420 343 -417
rect 356 -420 358 -417
rect 472 -420 474 -417
rect 497 -420 499 -417
rect 512 -420 514 -417
rect 549 -420 551 -417
rect 564 -420 566 -417
rect 65 -456 67 -453
rect 83 -456 85 -453
rect 110 -456 112 -453
rect 264 -459 266 -432
rect 264 -469 266 -466
rect 289 -485 291 -432
rect 304 -485 306 -432
rect 341 -485 343 -432
rect 356 -485 358 -432
rect 472 -459 474 -432
rect 472 -469 474 -466
rect 497 -485 499 -432
rect 512 -485 514 -432
rect 549 -485 551 -432
rect 564 -485 566 -432
rect 289 -494 291 -491
rect 304 -494 306 -491
rect 341 -494 343 -491
rect 356 -494 358 -491
rect 497 -494 499 -491
rect 512 -494 514 -491
rect 549 -494 551 -491
rect 564 -494 566 -491
rect -36 -499 -34 -496
rect -18 -499 -16 -496
rect 9 -499 11 -496
rect -759 -544 -757 -541
rect -744 -544 -742 -541
rect -707 -544 -705 -541
rect -692 -544 -690 -541
rect -551 -544 -549 -541
rect -536 -544 -534 -541
rect -499 -544 -497 -541
rect -484 -544 -482 -541
<< polycontact >>
rect -307 762 -302 766
rect -813 747 -808 751
rect -568 738 -563 742
rect -397 704 -392 708
rect -903 689 -898 693
rect -658 680 -653 684
rect -397 679 -393 683
rect -302 679 -297 683
rect -903 664 -899 668
rect -808 664 -803 668
rect -430 664 -426 668
rect -319 664 -314 668
rect -936 649 -932 653
rect -658 655 -654 659
rect -563 655 -558 659
rect -825 649 -820 653
rect -691 640 -687 644
rect -580 640 -575 644
rect -414 627 -410 631
rect -303 627 -299 631
rect -920 612 -916 616
rect -809 612 -805 616
rect -426 612 -422 616
rect -325 612 -321 616
rect -932 597 -928 601
rect -675 603 -671 607
rect -564 603 -560 607
rect -831 597 -827 601
rect -687 588 -683 592
rect -586 588 -582 592
rect -200 512 -196 517
rect -397 496 -392 500
rect -117 517 -113 522
rect -903 481 -898 485
rect -102 500 -98 505
rect -65 516 -61 520
rect -50 494 -46 498
rect 91 517 95 522
rect 106 500 110 505
rect 143 516 147 520
rect 158 494 162 498
rect -658 472 -653 476
rect -397 471 -393 475
rect -302 471 -297 475
rect -903 456 -899 460
rect -808 456 -803 460
rect -430 456 -426 460
rect -319 456 -314 460
rect -936 441 -932 445
rect -658 447 -654 451
rect -563 447 -558 451
rect -825 441 -820 445
rect -691 432 -687 436
rect -580 432 -575 436
rect -414 419 -410 423
rect -303 419 -299 423
rect -142 422 -138 427
rect -920 404 -916 408
rect -809 404 -805 408
rect -426 404 -422 408
rect -117 422 -113 426
rect -325 404 -321 408
rect -932 389 -928 393
rect -675 395 -671 399
rect -564 395 -560 399
rect -831 389 -827 393
rect -687 380 -683 384
rect -102 389 -98 393
rect -65 405 -61 409
rect -50 393 -46 397
rect 66 422 70 427
rect 91 422 95 426
rect 106 389 110 393
rect 143 405 147 409
rect 158 393 162 397
rect -586 380 -582 384
rect -931 300 -926 304
rect 74 307 78 312
rect -333 288 -329 292
rect -822 252 -818 257
rect -1021 242 -1016 246
rect -739 257 -735 262
rect -724 240 -720 245
rect -687 256 -683 260
rect -672 234 -668 238
rect -531 257 -527 262
rect -516 240 -512 245
rect -479 256 -475 260
rect -464 234 -460 238
rect -309 256 -305 260
rect -299 288 -295 292
rect -289 267 -285 271
rect -273 285 -269 289
rect 157 312 161 317
rect -255 288 -251 292
rect -173 269 -169 273
rect -148 229 -144 233
rect -1021 217 -1017 221
rect -926 217 -921 221
rect -136 267 -132 271
rect -122 255 -118 259
rect -103 267 -99 271
rect 172 295 176 300
rect 209 311 213 315
rect 224 289 228 293
rect 365 312 369 317
rect 380 295 384 300
rect 417 311 421 315
rect 432 289 436 293
rect -75 267 -71 271
rect -1054 202 -1050 206
rect 132 217 136 222
rect -943 202 -938 206
rect 157 217 161 221
rect -333 180 -329 184
rect -1038 165 -1034 169
rect -927 165 -923 169
rect -1050 150 -1046 154
rect -764 162 -760 167
rect -949 150 -945 154
rect -739 162 -735 166
rect -724 129 -720 133
rect -687 145 -683 149
rect -672 133 -668 137
rect -556 162 -552 167
rect -531 162 -527 166
rect -516 129 -512 133
rect -479 145 -475 149
rect -464 133 -460 137
rect -323 173 -319 177
rect -305 173 -301 177
rect 172 184 176 188
rect 209 200 213 204
rect 224 188 228 192
rect 340 217 344 222
rect 365 217 369 221
rect 380 184 384 188
rect 417 200 421 204
rect 432 188 436 192
rect -145 134 -141 138
rect -333 110 -329 114
rect -309 78 -305 82
rect -299 110 -295 114
rect -289 89 -285 93
rect -273 107 -269 111
rect -255 110 -251 114
rect -132 117 -128 121
rect -110 132 -106 136
rect -43 132 -38 137
rect -25 118 -20 123
rect 3 129 7 134
rect 66 103 70 107
rect -1021 34 -1016 38
rect -835 38 -831 43
rect -752 43 -748 48
rect -737 26 -733 31
rect -700 42 -696 46
rect -685 20 -681 24
rect -544 43 -540 48
rect -529 26 -525 31
rect -492 42 -488 46
rect -477 20 -473 24
rect 91 63 95 67
rect 103 101 107 105
rect 117 89 121 93
rect 136 101 140 105
rect 164 101 168 105
rect 295 80 299 85
rect 378 85 382 90
rect 393 68 397 73
rect 430 84 434 88
rect 445 62 449 66
rect 586 85 590 90
rect 601 68 605 73
rect 638 84 642 88
rect 653 62 657 66
rect -1021 9 -1017 13
rect -926 9 -921 13
rect -1054 -6 -1050 -2
rect -333 2 -329 6
rect -943 -6 -938 -2
rect -323 -5 -319 -1
rect -305 -5 -301 -1
rect -170 -8 -166 -4
rect -157 -25 -153 -21
rect -135 -10 -131 -6
rect -87 -22 -83 -18
rect -1038 -43 -1034 -39
rect -927 -43 -923 -39
rect -1050 -58 -1046 -54
rect -777 -52 -773 -47
rect -949 -58 -945 -54
rect -752 -52 -748 -48
rect -737 -85 -733 -81
rect -700 -69 -696 -65
rect -685 -81 -681 -77
rect -569 -52 -565 -47
rect -544 -52 -540 -48
rect -529 -85 -525 -81
rect -492 -69 -488 -65
rect -477 -81 -473 -77
rect -74 -39 -70 -35
rect -52 -24 -48 -20
rect 353 -10 357 -5
rect 378 -10 382 -6
rect 16 -55 21 -50
rect -333 -68 -329 -64
rect -309 -100 -305 -96
rect -299 -68 -295 -64
rect -289 -89 -285 -85
rect -273 -71 -269 -67
rect -255 -68 -251 -64
rect -179 -106 -175 -102
rect -166 -123 -162 -119
rect -144 -108 -140 -104
rect 34 -69 39 -64
rect 62 -58 66 -53
rect 126 -58 130 -54
rect 151 -98 155 -94
rect 163 -60 167 -56
rect 177 -72 181 -68
rect 196 -60 200 -56
rect 393 -43 397 -39
rect 430 -27 434 -23
rect 445 -39 449 -35
rect 561 -10 565 -5
rect 586 -10 590 -6
rect 601 -43 605 -39
rect 638 -27 642 -23
rect 653 -39 657 -35
rect 224 -60 228 -56
rect -85 -128 -80 -123
rect -837 -193 -833 -188
rect -754 -188 -750 -183
rect -739 -205 -735 -200
rect -702 -189 -698 -185
rect -687 -211 -683 -207
rect -546 -188 -542 -183
rect -531 -205 -527 -200
rect -494 -189 -490 -185
rect -479 -211 -475 -207
rect -67 -142 -62 -137
rect -39 -131 -35 -126
rect 289 -134 293 -129
rect 372 -129 376 -124
rect 387 -146 391 -141
rect 424 -130 428 -126
rect 439 -152 443 -148
rect 580 -129 584 -124
rect 595 -146 599 -141
rect 632 -130 636 -126
rect 647 -152 651 -148
rect -333 -176 -329 -172
rect -323 -183 -319 -179
rect -305 -183 -301 -179
rect -151 -225 -147 -221
rect -333 -246 -329 -242
rect -779 -283 -775 -278
rect -754 -283 -750 -279
rect -739 -316 -735 -312
rect -702 -300 -698 -296
rect -687 -312 -683 -308
rect -571 -283 -567 -278
rect -546 -283 -542 -279
rect -531 -316 -527 -312
rect -494 -300 -490 -296
rect -479 -312 -475 -308
rect -309 -278 -305 -274
rect -299 -246 -295 -242
rect -289 -267 -285 -263
rect -273 -249 -269 -245
rect -255 -246 -251 -242
rect -138 -242 -134 -238
rect -116 -227 -112 -223
rect -68 -239 -64 -235
rect -55 -256 -51 -252
rect -33 -241 -29 -237
rect 347 -224 351 -219
rect 15 -247 19 -243
rect 28 -264 32 -260
rect 50 -249 54 -245
rect 372 -224 376 -220
rect 387 -257 391 -253
rect 424 -241 428 -237
rect 439 -253 443 -249
rect 555 -224 559 -219
rect 580 -224 584 -220
rect 595 -257 599 -253
rect 632 -241 636 -237
rect 647 -253 651 -249
rect 96 -291 101 -286
rect -136 -341 -132 -337
rect -333 -354 -329 -350
rect -323 -361 -319 -357
rect -305 -361 -301 -357
rect -123 -358 -119 -354
rect -101 -343 -97 -339
rect 114 -305 119 -300
rect 142 -294 146 -289
rect -53 -355 -49 -351
rect -846 -408 -842 -403
rect -763 -403 -759 -398
rect -748 -420 -744 -415
rect -711 -404 -707 -400
rect -696 -426 -692 -422
rect -555 -403 -551 -398
rect -540 -420 -536 -415
rect -503 -404 -499 -400
rect -488 -426 -484 -422
rect -40 -372 -36 -368
rect -18 -357 -14 -353
rect 202 -358 206 -353
rect 285 -353 289 -348
rect 300 -370 304 -365
rect 337 -354 341 -350
rect 352 -376 356 -372
rect 493 -353 497 -348
rect 508 -370 512 -365
rect 545 -354 549 -350
rect 560 -376 564 -372
rect 60 -408 65 -403
rect -138 -435 -134 -431
rect -125 -452 -121 -448
rect -103 -437 -99 -433
rect -41 -451 -36 -446
rect -788 -498 -784 -493
rect -763 -498 -759 -494
rect -748 -531 -744 -527
rect -711 -515 -707 -511
rect -696 -527 -692 -523
rect -580 -498 -576 -493
rect -555 -498 -551 -494
rect -540 -531 -536 -527
rect -503 -515 -499 -511
rect -488 -527 -484 -523
rect -23 -465 -18 -460
rect 5 -454 9 -449
rect 78 -422 83 -417
rect 106 -411 110 -406
rect 260 -448 264 -443
rect 285 -448 289 -444
rect 300 -481 304 -477
rect 337 -465 341 -461
rect 352 -477 356 -473
rect 468 -448 472 -443
rect 493 -448 497 -444
rect 508 -481 512 -477
rect 545 -465 549 -461
rect 560 -477 564 -473
<< metal1 >>
rect -425 792 -302 796
rect -931 777 -808 781
rect -931 739 -927 777
rect -813 768 -808 777
rect -686 768 -563 772
rect -813 764 -682 768
rect -839 749 -831 753
rect -813 751 -808 764
rect -839 745 -836 749
rect -785 750 -772 754
rect -775 746 -772 750
rect -962 736 -927 739
rect -824 737 -797 741
rect -962 532 -958 736
rect -813 733 -809 737
rect -686 730 -682 764
rect -568 767 -563 768
rect -425 767 -421 792
rect -568 762 -421 767
rect -594 740 -586 744
rect -568 742 -563 762
rect -425 754 -421 762
rect -333 764 -325 768
rect -307 766 -302 792
rect -333 760 -330 764
rect -279 765 -266 769
rect -269 761 -266 765
rect -456 751 -421 754
rect -318 752 -291 756
rect -594 736 -591 740
rect -540 741 -527 745
rect -530 737 -527 741
rect -717 727 -682 730
rect -579 728 -552 732
rect -936 720 -831 723
rect -954 666 -946 670
rect -954 662 -950 666
rect -936 653 -932 720
rect -808 710 -803 718
rect -903 706 -803 710
rect -929 691 -921 695
rect -903 693 -898 706
rect -929 687 -926 691
rect -875 692 -862 696
rect -865 688 -862 692
rect -914 679 -887 683
rect -903 668 -899 679
rect -875 667 -862 671
rect -903 654 -887 658
rect -903 644 -899 654
rect -865 645 -862 667
rect -849 666 -841 670
rect -849 662 -845 666
rect -825 653 -821 672
rect -808 668 -803 706
rect -770 667 -757 671
rect -798 654 -782 658
rect -940 640 -899 644
rect -875 641 -862 645
rect -798 644 -794 654
rect -760 645 -757 667
rect -835 640 -794 644
rect -770 641 -757 645
rect -954 614 -946 618
rect -954 610 -950 614
rect -932 601 -928 640
rect -920 616 -916 623
rect -875 615 -862 619
rect -903 602 -887 606
rect -903 592 -899 602
rect -865 593 -862 615
rect -849 614 -841 618
rect -849 610 -845 614
rect -831 601 -827 640
rect -809 616 -805 622
rect -770 615 -757 619
rect -798 602 -782 606
rect -940 588 -899 592
rect -875 589 -862 593
rect -798 592 -794 602
rect -760 593 -757 615
rect -835 588 -794 592
rect -770 589 -757 593
rect -924 565 -920 588
rect -811 577 -807 588
rect -900 573 -807 577
rect -924 561 -820 565
rect -924 557 -920 561
rect -978 531 -958 532
rect -978 528 -821 531
rect -978 334 -971 528
rect -825 518 -821 528
rect -936 514 -821 518
rect -954 458 -946 462
rect -954 454 -950 458
rect -936 445 -932 514
rect -825 513 -821 514
rect -811 502 -807 573
rect -717 522 -713 727
rect -568 724 -564 728
rect -691 711 -586 714
rect -709 657 -701 661
rect -709 653 -705 657
rect -691 644 -687 711
rect -563 701 -558 709
rect -658 697 -558 701
rect -684 682 -676 686
rect -658 684 -653 697
rect -684 678 -681 682
rect -630 683 -617 687
rect -620 679 -617 683
rect -669 670 -642 674
rect -658 659 -654 670
rect -630 658 -617 662
rect -658 645 -642 649
rect -658 635 -654 645
rect -620 636 -617 658
rect -604 657 -596 661
rect -604 653 -600 657
rect -580 644 -576 663
rect -563 659 -558 697
rect -525 658 -512 662
rect -553 645 -537 649
rect -695 631 -654 635
rect -630 632 -617 636
rect -553 635 -549 645
rect -515 636 -512 658
rect -590 631 -549 635
rect -525 632 -512 636
rect -709 605 -701 609
rect -709 601 -705 605
rect -687 592 -683 631
rect -675 607 -671 614
rect -630 606 -617 610
rect -658 593 -642 597
rect -658 583 -654 593
rect -620 584 -617 606
rect -604 605 -596 609
rect -604 601 -600 605
rect -586 592 -582 631
rect -564 607 -560 613
rect -525 606 -512 610
rect -553 593 -537 597
rect -695 579 -654 583
rect -630 580 -617 584
rect -553 583 -549 593
rect -515 584 -512 606
rect -590 579 -549 583
rect -525 580 -512 584
rect -679 556 -675 579
rect -566 568 -562 579
rect -655 564 -562 568
rect -679 552 -575 556
rect -679 548 -675 552
rect -717 519 -576 522
rect -580 509 -576 519
rect -691 505 -576 509
rect -903 498 -803 502
rect -929 483 -921 487
rect -903 485 -898 498
rect -929 479 -926 483
rect -875 484 -862 488
rect -865 480 -862 484
rect -914 471 -887 475
rect -903 460 -899 471
rect -875 459 -862 463
rect -903 446 -887 450
rect -903 436 -899 446
rect -865 437 -862 459
rect -849 458 -841 462
rect -808 460 -803 498
rect -849 454 -845 458
rect -825 445 -821 460
rect -770 459 -757 463
rect -798 446 -782 450
rect -940 432 -899 436
rect -875 433 -862 437
rect -798 436 -794 446
rect -760 437 -757 459
rect -709 449 -701 453
rect -709 445 -705 449
rect -835 432 -794 436
rect -770 433 -757 437
rect -691 436 -687 505
rect -580 504 -576 505
rect -566 493 -562 564
rect -456 546 -452 751
rect -307 748 -303 752
rect -430 735 -325 738
rect -448 681 -440 685
rect -448 677 -444 681
rect -430 668 -426 735
rect -302 725 -297 733
rect -397 721 -297 725
rect -423 706 -415 710
rect -397 708 -392 721
rect -423 702 -420 706
rect -369 707 -356 711
rect -359 703 -356 707
rect -408 694 -381 698
rect -397 683 -393 694
rect -369 682 -356 686
rect -397 669 -381 673
rect -397 659 -393 669
rect -359 660 -356 682
rect -343 681 -335 685
rect -343 677 -339 681
rect -319 668 -315 687
rect -302 683 -297 721
rect -264 682 -251 686
rect -292 669 -276 673
rect -434 655 -393 659
rect -369 656 -356 660
rect -292 659 -288 669
rect -254 660 -251 682
rect -329 655 -288 659
rect -264 656 -251 660
rect -448 629 -440 633
rect -448 625 -444 629
rect -426 616 -422 655
rect -414 631 -410 638
rect -369 630 -356 634
rect -397 617 -381 621
rect -397 607 -393 617
rect -359 608 -356 630
rect -343 629 -335 633
rect -343 625 -339 629
rect -325 616 -321 655
rect -303 631 -299 637
rect -264 630 -251 634
rect -292 617 -276 621
rect -434 603 -393 607
rect -369 604 -356 608
rect -292 607 -288 617
rect -254 608 -251 630
rect -329 603 -288 607
rect -264 604 -251 608
rect -418 580 -414 603
rect -305 592 -301 603
rect -394 588 -301 592
rect -418 576 -314 580
rect -418 572 -414 576
rect -456 543 -315 546
rect -319 533 -315 543
rect -430 529 -315 533
rect -658 489 -558 493
rect -684 474 -676 478
rect -658 476 -653 489
rect -684 470 -681 474
rect -630 475 -617 479
rect -620 471 -617 475
rect -669 462 -642 466
rect -658 451 -654 462
rect -630 450 -617 454
rect -658 437 -642 441
rect -954 406 -946 410
rect -954 402 -950 406
rect -932 393 -928 432
rect -920 408 -916 415
rect -875 407 -862 411
rect -903 394 -887 398
rect -903 384 -899 394
rect -865 385 -862 407
rect -849 406 -841 410
rect -849 402 -845 406
rect -831 393 -827 432
rect -658 427 -654 437
rect -620 428 -617 450
rect -604 449 -596 453
rect -563 451 -558 489
rect -448 473 -440 477
rect -448 469 -444 473
rect -430 460 -426 529
rect -319 528 -315 529
rect -305 517 -301 588
rect -120 565 -90 568
rect -120 555 -116 565
rect -94 555 -90 565
rect -203 550 -195 553
rect -203 540 -199 550
rect -68 565 -38 568
rect -68 555 -64 565
rect -42 555 -38 565
rect 88 565 118 568
rect 88 555 92 565
rect 114 555 118 565
rect 140 565 170 568
rect 140 555 144 565
rect 166 555 170 565
rect -397 513 -297 517
rect -423 498 -415 502
rect -397 500 -392 513
rect -423 494 -420 498
rect -369 499 -356 503
rect -359 495 -356 499
rect -408 486 -381 490
rect -397 475 -393 486
rect -369 474 -356 478
rect -397 461 -381 465
rect -604 445 -600 449
rect -580 436 -576 451
rect -525 450 -512 454
rect -397 451 -393 461
rect -359 452 -356 474
rect -343 473 -335 477
rect -302 475 -297 513
rect -230 512 -200 517
rect -190 516 -186 528
rect -107 531 -103 543
rect -55 531 -51 543
rect 101 531 105 543
rect 153 531 157 543
rect -107 527 -89 531
rect -55 527 -37 531
rect 101 527 119 531
rect 153 527 171 531
rect -159 517 -117 522
rect -190 512 -182 516
rect -343 469 -339 473
rect -319 460 -315 475
rect -264 474 -251 478
rect -292 461 -276 465
rect -553 437 -537 441
rect -695 423 -654 427
rect -630 424 -617 428
rect -553 427 -549 437
rect -515 428 -512 450
rect -434 447 -393 451
rect -369 448 -356 452
rect -292 451 -288 461
rect -254 452 -251 474
rect -329 447 -288 451
rect -264 448 -251 452
rect -590 423 -549 427
rect -525 424 -512 428
rect -809 408 -805 414
rect -770 407 -757 411
rect -798 394 -782 398
rect -940 380 -899 384
rect -875 381 -862 385
rect -798 384 -794 394
rect -760 385 -757 407
rect -709 397 -701 401
rect -709 393 -705 397
rect -835 380 -794 384
rect -770 381 -757 385
rect -687 384 -683 423
rect -675 399 -671 406
rect -630 398 -617 402
rect -658 385 -642 389
rect -924 357 -920 380
rect -811 369 -807 380
rect -658 375 -654 385
rect -620 376 -617 398
rect -604 397 -596 401
rect -604 393 -600 397
rect -586 384 -582 423
rect -448 421 -440 425
rect -448 417 -444 421
rect -426 408 -422 447
rect -414 423 -410 430
rect -369 422 -356 426
rect -564 399 -560 405
rect -397 409 -381 413
rect -525 398 -512 402
rect -397 399 -393 409
rect -359 400 -356 422
rect -343 421 -335 425
rect -343 417 -339 421
rect -325 408 -321 447
rect -303 423 -299 429
rect -264 422 -251 426
rect -292 409 -276 413
rect -553 385 -537 389
rect -695 371 -654 375
rect -630 372 -617 376
rect -553 375 -549 385
rect -515 376 -512 398
rect -434 395 -393 399
rect -369 396 -356 400
rect -292 399 -288 409
rect -254 400 -251 422
rect -329 395 -288 399
rect -264 396 -251 400
rect -230 398 -226 512
rect -190 501 -186 512
rect -202 489 -198 494
rect -202 486 -194 489
rect -590 371 -549 375
rect -525 372 -512 376
rect -418 372 -414 395
rect -305 384 -301 395
rect -230 394 -185 398
rect -394 380 -301 384
rect -900 367 -807 369
rect -900 366 -733 367
rect -900 365 -732 366
rect -811 362 -732 365
rect -924 353 -820 357
rect -924 349 -920 353
rect -1049 331 -926 334
rect -1049 330 -847 331
rect -1049 292 -1045 330
rect -931 326 -847 330
rect -957 302 -949 306
rect -931 304 -926 326
rect -957 298 -954 302
rect -903 303 -890 307
rect -893 299 -890 303
rect -1080 289 -1045 292
rect -942 290 -915 294
rect -1080 84 -1076 289
rect -931 286 -927 290
rect -1054 273 -949 276
rect -1072 219 -1064 223
rect -1072 215 -1068 219
rect -1054 206 -1050 273
rect -926 263 -921 271
rect -1021 259 -921 263
rect -1047 244 -1039 248
rect -1021 246 -1016 259
rect -1047 240 -1044 244
rect -993 245 -980 249
rect -983 241 -980 245
rect -1032 232 -1005 236
rect -1021 221 -1017 232
rect -993 220 -980 224
rect -1021 207 -1005 211
rect -1021 197 -1017 207
rect -983 198 -980 220
rect -967 219 -959 223
rect -967 215 -963 219
rect -943 206 -939 225
rect -926 221 -921 259
rect -853 257 -847 326
rect -736 328 -732 362
rect -679 348 -675 371
rect -566 360 -562 371
rect -418 368 -314 372
rect -418 364 -414 368
rect -655 356 -562 360
rect -566 352 -369 356
rect -305 354 -301 380
rect -188 367 -185 394
rect -172 393 -169 494
rect -159 465 -155 517
rect -121 500 -102 504
rect -93 498 -89 527
rect -71 516 -65 520
rect -41 518 -37 527
rect 49 518 91 522
rect -41 517 91 518
rect -41 514 53 517
rect -93 494 -50 498
rect -93 490 -89 494
rect -41 490 -37 514
rect -119 480 -115 484
rect -67 480 -63 484
rect -119 476 -111 480
rect -67 476 -59 480
rect -158 460 -155 465
rect -159 427 -155 460
rect -145 460 -137 463
rect -120 460 -90 463
rect -145 450 -141 460
rect -120 450 -116 460
rect -94 450 -90 460
rect -68 460 -38 463
rect -68 450 -64 460
rect -42 450 -38 460
rect -159 422 -142 427
rect -132 426 -128 438
rect -107 426 -103 438
rect -55 426 -51 438
rect -132 422 -117 426
rect -107 422 -89 426
rect -55 422 -37 426
rect -132 411 -128 422
rect -144 399 -140 404
rect -144 396 -136 399
rect -93 397 -89 422
rect -72 405 -65 409
rect -41 405 -37 422
rect -26 425 -22 514
rect -14 405 -10 505
rect 20 500 38 504
rect -41 401 -6 405
rect -93 393 -50 397
rect -172 389 -102 393
rect -93 385 -89 393
rect -41 385 -37 401
rect -119 375 -115 379
rect -67 375 -63 379
rect -119 371 -111 375
rect -67 371 -59 375
rect 20 367 23 500
rect 33 393 37 500
rect 49 427 53 514
rect 91 500 106 504
rect 115 498 119 527
rect 137 516 143 520
rect 167 518 171 527
rect 167 514 205 518
rect 115 494 158 498
rect 115 490 119 494
rect 167 490 171 514
rect 89 480 93 484
rect 141 480 145 484
rect 89 476 97 480
rect 141 476 149 480
rect 63 460 71 463
rect 88 460 118 463
rect 63 450 67 460
rect 88 450 92 460
rect 114 450 118 460
rect 140 460 170 463
rect 140 450 144 460
rect 166 450 170 460
rect 49 422 66 427
rect 76 426 80 438
rect 101 426 105 438
rect 153 426 157 438
rect 76 422 91 426
rect 101 422 119 426
rect 153 422 171 426
rect 76 411 80 422
rect 64 399 68 404
rect 64 396 72 399
rect 115 397 119 422
rect 136 405 143 409
rect 167 405 171 422
rect 182 425 186 514
rect 194 405 198 505
rect 167 401 202 405
rect 115 393 158 397
rect 33 389 106 393
rect -188 363 23 367
rect -679 344 -575 348
rect -679 340 -675 344
rect -373 347 -369 352
rect -359 351 -301 354
rect -736 324 -380 328
rect -742 305 -712 308
rect -742 295 -738 305
rect -716 295 -712 305
rect -825 290 -817 293
rect -825 280 -821 290
rect -690 305 -660 308
rect -690 295 -686 305
rect -664 295 -660 305
rect -534 305 -504 308
rect -534 295 -530 305
rect -508 295 -504 305
rect -482 305 -452 308
rect -482 295 -478 305
rect -456 295 -452 305
rect -853 255 -822 257
rect -852 252 -822 255
rect -812 256 -808 268
rect -729 271 -725 283
rect -677 271 -673 283
rect -521 271 -517 283
rect -469 271 -465 283
rect -729 267 -711 271
rect -677 267 -659 271
rect -521 267 -503 271
rect -469 267 -451 271
rect -789 257 -739 262
rect -812 252 -804 256
rect -888 220 -875 224
rect -916 207 -900 211
rect -1058 193 -1017 197
rect -993 194 -980 198
rect -916 197 -912 207
rect -878 198 -875 220
rect -953 193 -912 197
rect -888 194 -875 198
rect -1072 167 -1064 171
rect -1072 163 -1068 167
rect -1050 154 -1046 193
rect -1038 169 -1034 176
rect -993 168 -980 172
rect -1021 155 -1005 159
rect -1021 145 -1017 155
rect -983 146 -980 168
rect -967 167 -959 171
rect -967 163 -963 167
rect -949 154 -945 193
rect -927 169 -923 175
rect -888 168 -875 172
rect -916 155 -900 159
rect -1058 141 -1017 145
rect -993 142 -980 146
rect -916 145 -912 155
rect -878 146 -875 168
rect -953 141 -912 145
rect -888 142 -875 146
rect -1042 118 -1038 141
rect -929 130 -925 141
rect -1018 126 -925 130
rect -1042 114 -938 118
rect -1042 110 -1038 114
rect -1080 81 -939 84
rect -1080 -138 -1076 81
rect -943 71 -939 81
rect -1054 67 -939 71
rect -1072 11 -1064 15
rect -1072 7 -1068 11
rect -1054 -2 -1050 67
rect -943 66 -939 67
rect -929 55 -925 126
rect -852 139 -848 252
rect -812 241 -808 252
rect -824 229 -820 234
rect -824 226 -816 229
rect -852 138 -847 139
rect -852 134 -807 138
rect -1021 51 -921 55
rect -1047 36 -1039 40
rect -1021 38 -1016 51
rect -1047 32 -1044 36
rect -993 37 -980 41
rect -983 33 -980 37
rect -1032 24 -1005 28
rect -1021 13 -1017 24
rect -993 12 -980 16
rect -1021 -1 -1005 3
rect -1021 -11 -1017 -1
rect -983 -10 -980 12
rect -967 11 -959 15
rect -926 13 -921 51
rect -852 43 -847 134
rect -810 107 -807 134
rect -794 133 -791 234
rect -781 167 -777 257
rect -743 240 -724 244
rect -715 238 -711 267
rect -693 256 -687 260
rect -663 258 -659 267
rect -573 258 -531 262
rect -663 257 -531 258
rect -663 254 -569 257
rect -715 234 -672 238
rect -715 230 -711 234
rect -663 230 -659 254
rect -741 220 -737 224
rect -689 220 -685 224
rect -741 216 -733 220
rect -689 216 -681 220
rect -767 200 -759 203
rect -742 200 -712 203
rect -767 190 -763 200
rect -742 190 -738 200
rect -716 190 -712 200
rect -690 200 -660 203
rect -690 190 -686 200
rect -664 190 -660 200
rect -781 162 -764 167
rect -754 166 -750 178
rect -729 166 -725 178
rect -677 166 -673 178
rect -754 162 -739 166
rect -729 162 -711 166
rect -677 162 -659 166
rect -754 151 -750 162
rect -766 139 -762 144
rect -766 136 -758 139
rect -715 137 -711 162
rect -694 145 -687 149
rect -663 145 -659 162
rect -648 165 -644 254
rect -636 145 -632 245
rect -602 240 -584 244
rect -663 141 -628 145
rect -715 133 -672 137
rect -794 129 -724 133
rect -715 125 -711 133
rect -663 125 -659 141
rect -741 115 -737 119
rect -689 115 -685 119
rect -741 111 -733 115
rect -689 111 -681 115
rect -602 107 -599 240
rect -589 133 -585 240
rect -573 167 -569 254
rect -531 240 -516 244
rect -507 238 -503 267
rect -485 256 -479 260
rect -455 258 -451 267
rect -455 254 -391 258
rect -507 234 -464 238
rect -507 230 -503 234
rect -455 230 -451 254
rect -533 220 -529 224
rect -481 220 -477 224
rect -533 216 -525 220
rect -481 216 -473 220
rect -559 200 -551 203
rect -534 200 -504 203
rect -559 190 -555 200
rect -534 190 -530 200
rect -508 190 -504 200
rect -482 200 -452 203
rect -482 190 -478 200
rect -456 190 -452 200
rect -573 162 -556 167
rect -546 166 -542 178
rect -521 166 -517 178
rect -469 166 -465 178
rect -546 162 -531 166
rect -521 162 -503 166
rect -469 162 -451 166
rect -546 151 -542 162
rect -558 139 -554 144
rect -558 136 -550 139
rect -507 137 -503 162
rect -486 145 -479 149
rect -455 145 -451 162
rect -440 165 -436 254
rect -428 145 -424 245
rect -455 141 -420 145
rect -507 133 -464 137
rect -589 129 -516 133
rect -507 125 -503 133
rect -455 125 -451 141
rect -533 115 -529 119
rect -481 115 -477 119
rect -395 115 -391 254
rect -533 111 -525 115
rect -481 111 -473 115
rect -384 114 -380 324
rect -359 292 -355 351
rect -341 321 -243 325
rect -335 318 -331 321
rect -311 318 -307 321
rect -271 318 -267 321
rect -253 318 -249 321
rect 47 312 50 389
rect 115 385 119 393
rect 167 385 171 401
rect 89 375 93 379
rect 141 375 145 379
rect 89 371 97 375
rect 141 371 149 375
rect 154 360 184 363
rect 154 350 158 360
rect 180 350 184 360
rect 71 345 79 348
rect 71 335 75 345
rect 206 360 236 363
rect 206 350 210 360
rect 232 350 236 360
rect 362 360 392 363
rect 362 350 366 360
rect 388 350 392 360
rect 414 360 444 363
rect 414 350 418 360
rect 440 350 444 360
rect -183 305 -163 309
rect -152 305 -94 309
rect -81 305 -61 309
rect 44 307 74 312
rect 84 311 88 323
rect 167 326 171 338
rect 219 326 223 338
rect 375 326 379 338
rect 427 326 431 338
rect 167 322 185 326
rect 219 322 237 326
rect 375 322 393 326
rect 427 322 445 326
rect 115 312 157 317
rect 84 307 92 311
rect -325 292 -321 298
rect -291 292 -287 298
rect -359 288 -333 292
rect -325 288 -299 292
rect -291 288 -277 292
rect -263 289 -259 298
rect -176 296 -172 305
rect -151 296 -147 305
rect -98 296 -94 305
rect -72 296 -68 305
rect -355 177 -351 288
rect -341 266 -338 288
rect -325 285 -321 288
rect -335 272 -331 275
rect -335 269 -321 272
rect -312 267 -289 271
rect -312 266 -308 267
rect -341 263 -308 266
rect -281 264 -277 288
rect -269 285 -259 289
rect -251 288 -243 292
rect -253 272 -249 275
rect -262 268 -249 272
rect -301 260 -258 264
rect -343 256 -309 260
rect -348 184 -344 255
rect -322 223 -319 256
rect -301 250 -297 260
rect -291 253 -267 257
rect -291 250 -287 253
rect -271 250 -267 253
rect -311 237 -307 240
rect -291 237 -287 240
rect -311 233 -287 237
rect -281 230 -277 240
rect -313 226 -266 230
rect -246 223 -243 288
rect -214 269 -173 273
rect -164 271 -160 289
rect -126 272 -122 289
rect -322 220 -243 223
rect -236 254 -194 258
rect -341 213 -287 217
rect -335 210 -331 213
rect -315 210 -311 213
rect -307 210 -303 213
rect -325 184 -321 190
rect -348 180 -333 184
rect -325 180 -311 184
rect -315 177 -311 180
rect -297 177 -293 190
rect -236 177 -232 254
rect -198 233 -194 254
rect -187 241 -183 269
rect -164 267 -136 271
rect -126 268 -109 272
rect -84 271 -80 289
rect -164 259 -160 267
rect -150 255 -122 259
rect -176 247 -172 250
rect -176 244 -165 247
rect -150 241 -146 255
rect -187 238 -146 241
rect -113 239 -109 268
rect -99 267 -80 271
rect -71 267 -59 271
rect -84 260 -80 267
rect -72 248 -68 251
rect -76 244 -68 248
rect -139 235 -98 239
rect -198 229 -148 233
rect -162 195 -158 229
rect -139 223 -135 235
rect -127 227 -95 232
rect -127 223 -122 227
rect -100 223 -95 227
rect -152 208 -147 213
rect -127 208 -122 213
rect -152 204 -122 208
rect -113 202 -109 213
rect -119 198 -109 202
rect -63 196 -59 267
rect -77 195 -59 196
rect -162 191 -59 195
rect 44 193 48 307
rect 84 296 88 307
rect 72 284 76 289
rect 72 281 80 284
rect 44 189 89 193
rect -355 173 -323 177
rect -315 173 -305 177
rect -297 173 -232 177
rect -315 170 -311 173
rect -297 170 -293 173
rect -335 157 -331 160
rect -307 157 -303 160
rect -341 153 -287 157
rect -341 143 -243 147
rect -335 140 -331 143
rect -311 140 -307 143
rect -271 140 -267 143
rect -253 140 -249 143
rect -236 138 -232 173
rect -148 169 -110 174
rect -148 160 -143 169
rect -124 160 -120 169
rect -114 160 -110 169
rect -48 169 4 173
rect -133 140 -129 149
rect -236 137 -145 138
rect -236 135 -203 137
rect -198 135 -145 137
rect -133 136 -121 140
rect -102 136 -98 149
rect -48 159 -42 169
rect -1 159 4 169
rect 86 162 89 189
rect 102 188 105 289
rect 115 222 119 312
rect 153 295 172 299
rect 181 293 185 322
rect 203 311 209 315
rect 233 313 237 322
rect 323 313 365 317
rect 233 312 365 313
rect 233 309 327 312
rect 181 289 224 293
rect 181 285 185 289
rect 233 285 237 309
rect 155 275 159 279
rect 207 275 211 279
rect 155 271 163 275
rect 207 271 215 275
rect 129 255 137 258
rect 154 255 184 258
rect 129 245 133 255
rect 154 245 158 255
rect 180 245 184 255
rect 206 255 236 258
rect 206 245 210 255
rect 232 245 236 255
rect 115 217 132 222
rect 142 221 146 233
rect 167 221 171 233
rect 219 221 223 233
rect 142 217 157 221
rect 167 217 185 221
rect 219 217 237 221
rect 142 206 146 217
rect 130 194 134 199
rect 130 191 138 194
rect 181 192 185 217
rect 202 200 209 204
rect 233 200 237 217
rect 248 220 252 309
rect 260 200 264 300
rect 294 295 312 299
rect 233 196 268 200
rect 181 188 224 192
rect 102 184 172 188
rect 181 180 185 188
rect 233 180 237 196
rect 155 170 159 174
rect 207 170 211 174
rect 155 166 163 170
rect 207 166 215 170
rect 294 162 297 295
rect 307 188 311 295
rect 323 222 327 309
rect 365 295 380 299
rect 389 293 393 322
rect 411 311 417 315
rect 441 313 445 322
rect 441 309 478 313
rect 389 289 432 293
rect 389 285 393 289
rect 441 285 445 309
rect 363 275 367 279
rect 415 275 419 279
rect 363 271 371 275
rect 415 271 423 275
rect 337 255 345 258
rect 362 255 392 258
rect 337 245 341 255
rect 362 245 366 255
rect 388 245 392 255
rect 414 255 444 258
rect 414 245 418 255
rect 440 245 444 255
rect 323 217 340 222
rect 350 221 354 233
rect 375 221 379 233
rect 427 221 431 233
rect 350 217 365 221
rect 375 217 393 221
rect 427 217 445 221
rect 350 206 354 217
rect 338 194 342 199
rect 338 191 346 194
rect 389 192 393 217
rect 410 200 417 204
rect 441 200 445 217
rect 456 220 460 309
rect 468 200 472 300
rect 441 196 476 200
rect 389 188 432 192
rect 307 184 380 188
rect 389 180 393 188
rect 441 180 445 196
rect 363 170 367 174
rect 415 170 419 174
rect 363 166 371 170
rect 415 166 423 170
rect 86 158 297 162
rect -125 132 -110 136
rect -102 132 -43 136
rect -14 134 -9 148
rect -236 120 -224 121
rect -219 120 -132 121
rect -325 114 -321 120
rect -291 114 -287 120
rect -384 110 -333 114
rect -325 110 -299 114
rect -291 110 -277 114
rect -263 111 -259 120
rect -236 117 -132 120
rect -810 103 -599 107
rect -755 91 -725 94
rect -755 81 -751 91
rect -729 81 -725 91
rect -838 76 -830 79
rect -838 66 -834 76
rect -703 91 -673 94
rect -703 81 -699 91
rect -677 81 -673 91
rect -547 91 -517 94
rect -547 81 -543 91
rect -521 81 -517 91
rect -495 91 -465 94
rect -495 81 -491 91
rect -469 81 -465 91
rect -865 38 -835 43
rect -825 42 -821 54
rect -742 57 -738 69
rect -690 57 -686 69
rect -534 57 -530 69
rect -482 57 -478 69
rect -742 53 -724 57
rect -690 53 -672 57
rect -534 53 -516 57
rect -482 53 -464 57
rect -802 43 -752 48
rect -825 38 -817 42
rect -967 7 -963 11
rect -943 -2 -939 13
rect -888 12 -875 16
rect -916 -1 -900 3
rect -1058 -15 -1017 -11
rect -993 -14 -980 -10
rect -916 -11 -912 -1
rect -878 -10 -875 12
rect -953 -15 -912 -11
rect -888 -14 -875 -10
rect -1072 -41 -1064 -37
rect -1072 -45 -1068 -41
rect -1050 -54 -1046 -15
rect -1038 -39 -1034 -32
rect -993 -40 -980 -36
rect -1021 -53 -1005 -49
rect -1021 -63 -1017 -53
rect -983 -62 -980 -40
rect -967 -41 -959 -37
rect -967 -45 -963 -41
rect -949 -54 -945 -15
rect -927 -39 -923 -33
rect -888 -40 -875 -36
rect -916 -53 -900 -49
rect -1058 -67 -1017 -63
rect -993 -66 -980 -62
rect -916 -63 -912 -53
rect -878 -62 -875 -40
rect -953 -67 -912 -63
rect -888 -66 -875 -62
rect -1042 -90 -1038 -67
rect -929 -78 -925 -67
rect -1018 -82 -925 -78
rect -865 -76 -861 38
rect -825 27 -821 38
rect -837 15 -833 20
rect -837 12 -829 15
rect -865 -80 -820 -76
rect -1042 -94 -938 -90
rect -1042 -98 -1038 -94
rect -929 -115 -925 -82
rect -823 -107 -820 -80
rect -807 -81 -804 20
rect -794 -47 -790 43
rect -756 26 -737 30
rect -728 24 -724 53
rect -706 42 -700 46
rect -676 44 -672 53
rect -586 44 -544 48
rect -676 43 -544 44
rect -676 40 -582 43
rect -728 20 -685 24
rect -728 16 -724 20
rect -676 16 -672 40
rect -754 6 -750 10
rect -702 6 -698 10
rect -754 2 -746 6
rect -702 2 -694 6
rect -780 -14 -772 -11
rect -755 -14 -725 -11
rect -780 -24 -776 -14
rect -755 -24 -751 -14
rect -729 -24 -725 -14
rect -703 -14 -673 -11
rect -703 -24 -699 -14
rect -677 -24 -673 -14
rect -794 -52 -777 -47
rect -767 -48 -763 -36
rect -742 -48 -738 -36
rect -690 -48 -686 -36
rect -767 -52 -752 -48
rect -742 -52 -724 -48
rect -690 -52 -672 -48
rect -767 -63 -763 -52
rect -779 -75 -775 -70
rect -779 -78 -771 -75
rect -728 -77 -724 -52
rect -707 -69 -700 -65
rect -676 -69 -672 -52
rect -661 -49 -657 40
rect -649 -69 -645 31
rect -615 26 -597 30
rect -676 -73 -641 -69
rect -728 -81 -685 -77
rect -807 -85 -737 -81
rect -728 -89 -724 -81
rect -676 -89 -672 -73
rect -754 -99 -750 -95
rect -702 -99 -698 -95
rect -754 -103 -746 -99
rect -702 -103 -694 -99
rect -615 -107 -612 26
rect -602 -81 -598 26
rect -586 -47 -582 40
rect -544 26 -529 30
rect -520 24 -516 53
rect -498 42 -492 46
rect -468 44 -464 53
rect -468 40 -362 44
rect -520 20 -477 24
rect -520 16 -516 20
rect -468 16 -464 40
rect -546 6 -542 10
rect -494 6 -490 10
rect -546 2 -538 6
rect -494 2 -486 6
rect -572 -14 -564 -11
rect -547 -14 -517 -11
rect -572 -24 -568 -14
rect -547 -24 -543 -14
rect -521 -24 -517 -14
rect -495 -14 -465 -11
rect -495 -24 -491 -14
rect -469 -24 -465 -14
rect -586 -52 -569 -47
rect -559 -48 -555 -36
rect -534 -48 -530 -36
rect -482 -48 -478 -36
rect -559 -52 -544 -48
rect -534 -52 -516 -48
rect -482 -52 -464 -48
rect -559 -63 -555 -52
rect -571 -75 -567 -70
rect -571 -78 -563 -75
rect -520 -77 -516 -52
rect -499 -69 -492 -65
rect -468 -69 -464 -52
rect -453 -49 -449 40
rect -441 -69 -437 31
rect -365 -65 -362 40
rect -355 -1 -351 110
rect -341 88 -338 110
rect -325 107 -321 110
rect -335 94 -331 97
rect -335 91 -321 94
rect -312 89 -289 93
rect -312 88 -308 89
rect -341 85 -308 88
rect -281 86 -277 110
rect -269 107 -259 111
rect -251 110 -243 114
rect -253 94 -249 97
rect -262 90 -249 94
rect -301 82 -258 86
rect -343 78 -309 82
rect -348 6 -344 77
rect -322 45 -319 78
rect -301 72 -297 82
rect -291 75 -267 79
rect -291 72 -287 75
rect -271 72 -267 75
rect -311 59 -307 62
rect -291 59 -287 62
rect -311 55 -287 59
rect -281 52 -277 62
rect -313 48 -266 52
rect -246 45 -243 110
rect -236 87 -233 117
rect -125 108 -121 132
rect -102 109 -98 132
rect -14 129 3 134
rect -66 118 -25 122
rect -147 95 -143 100
rect -111 95 -107 101
rect -147 91 -107 95
rect -66 67 -62 118
rect -14 103 -9 129
rect -30 98 -9 103
rect 12 126 16 148
rect 56 139 76 143
rect 87 139 145 143
rect 158 139 178 143
rect 63 130 67 139
rect 88 130 92 139
rect 141 130 145 139
rect 167 130 171 139
rect 12 121 42 126
rect -30 95 -25 98
rect 12 95 16 121
rect 38 107 42 121
rect 38 103 66 107
rect 75 105 79 123
rect 113 106 117 123
rect -45 79 -40 87
rect -14 79 -9 87
rect 1 79 6 87
rect -45 74 6 79
rect 52 75 56 103
rect 75 101 103 105
rect 113 102 130 106
rect 155 105 159 123
rect 75 93 79 101
rect 89 89 117 93
rect 63 81 67 84
rect 63 78 74 81
rect 89 75 93 89
rect 52 72 93 75
rect 126 73 130 102
rect 140 101 159 105
rect 168 101 180 105
rect 155 94 159 101
rect 167 82 171 85
rect 163 78 171 82
rect 100 69 141 73
rect -322 42 -243 45
rect -233 62 -62 67
rect 53 63 91 67
rect -341 35 -287 39
rect -335 32 -331 35
rect -315 32 -311 35
rect -307 32 -303 35
rect -325 6 -321 12
rect -348 2 -333 6
rect -325 2 -311 6
rect -315 -1 -311 2
rect -297 -1 -293 12
rect -233 -1 -229 62
rect 53 46 57 63
rect -93 41 57 46
rect -203 -1 -199 32
rect -173 27 -135 32
rect -173 18 -168 27
rect -149 18 -145 27
rect -139 18 -135 27
rect 77 29 81 63
rect 100 57 104 69
rect 112 61 144 66
rect 112 57 117 61
rect 139 57 144 61
rect 87 42 92 47
rect 112 42 117 47
rect 87 38 117 42
rect 126 36 130 47
rect 120 32 130 36
rect 176 30 180 101
rect 272 85 275 158
rect 375 133 405 136
rect 375 123 379 133
rect 401 123 405 133
rect 292 118 300 121
rect 292 108 296 118
rect 427 133 457 136
rect 427 123 431 133
rect 453 123 457 133
rect 583 133 613 136
rect 583 123 587 133
rect 609 123 613 133
rect 635 133 665 136
rect 635 123 639 133
rect 661 123 665 133
rect 162 29 180 30
rect 77 25 180 29
rect 265 80 295 85
rect 305 84 309 96
rect 388 99 392 111
rect 440 99 444 111
rect 596 99 600 111
rect 648 99 652 111
rect 388 95 406 99
rect 440 95 458 99
rect 596 95 614 99
rect 648 95 666 99
rect 336 85 378 90
rect 305 80 313 84
rect -355 -5 -323 -1
rect -315 -5 -305 -1
rect -297 -5 -229 -1
rect -315 -8 -311 -5
rect -297 -8 -293 -5
rect -335 -21 -331 -18
rect -307 -21 -303 -18
rect -341 -25 -282 -21
rect -233 -30 -229 -5
rect -215 -4 -199 -1
rect -158 -2 -154 7
rect -215 -5 -170 -4
rect -341 -35 -243 -31
rect -335 -38 -331 -35
rect -311 -38 -307 -35
rect -271 -38 -267 -35
rect -253 -38 -249 -35
rect -215 -46 -212 -5
rect -203 -8 -170 -5
rect -158 -6 -146 -2
rect -150 -10 -135 -6
rect -127 -8 -123 7
rect -90 13 -52 18
rect -90 4 -85 13
rect -66 4 -62 13
rect -56 4 -52 13
rect -173 -21 -160 -20
rect -173 -24 -157 -21
rect -162 -25 -157 -24
rect -150 -34 -146 -10
rect -127 -12 -105 -8
rect -127 -33 -123 -12
rect -108 -18 -105 -12
rect -75 -16 -71 -7
rect -108 -21 -87 -18
rect -75 -20 -63 -16
rect -67 -24 -52 -20
rect -44 -22 -40 -7
rect 11 -18 63 -14
rect -103 -39 -74 -36
rect -172 -47 -168 -42
rect -136 -47 -132 -41
rect -172 -51 -132 -47
rect -325 -64 -321 -58
rect -291 -64 -287 -58
rect -359 -65 -333 -64
rect -365 -68 -333 -65
rect -325 -68 -299 -64
rect -291 -68 -277 -64
rect -263 -67 -259 -58
rect -103 -59 -100 -39
rect -67 -48 -63 -24
rect -44 -26 -7 -22
rect -44 -47 -40 -26
rect -239 -62 -100 -59
rect -11 -50 -7 -26
rect 11 -28 17 -18
rect 58 -28 63 -18
rect 116 -22 136 -18
rect 147 -22 205 -18
rect 218 -22 238 -18
rect 123 -31 127 -22
rect 148 -31 152 -22
rect 201 -31 205 -22
rect 227 -31 231 -22
rect 265 -34 269 80
rect 305 69 309 80
rect 293 57 297 62
rect 293 54 301 57
rect 265 -38 310 -34
rect -11 -54 16 -50
rect 45 -53 50 -39
rect -89 -61 -85 -56
rect -53 -61 -49 -55
rect -468 -73 -433 -69
rect -520 -81 -477 -77
rect -602 -85 -529 -81
rect -520 -89 -516 -81
rect -468 -89 -464 -73
rect -546 -99 -542 -95
rect -494 -99 -490 -95
rect -546 -103 -538 -99
rect -494 -103 -486 -99
rect -823 -111 -612 -107
rect -929 -118 -415 -115
rect -1080 -142 -863 -138
rect -1080 -143 -886 -142
rect -867 -188 -863 -142
rect -757 -140 -727 -137
rect -757 -150 -753 -140
rect -731 -150 -727 -140
rect -840 -155 -832 -152
rect -840 -165 -836 -155
rect -705 -140 -675 -137
rect -705 -150 -701 -140
rect -679 -150 -675 -140
rect -549 -140 -519 -137
rect -549 -150 -545 -140
rect -523 -150 -519 -140
rect -497 -140 -467 -137
rect -497 -150 -493 -140
rect -471 -150 -467 -140
rect -867 -193 -837 -188
rect -827 -189 -823 -177
rect -744 -174 -740 -162
rect -692 -174 -688 -162
rect -536 -174 -532 -162
rect -484 -174 -480 -162
rect -744 -178 -726 -174
rect -692 -178 -674 -174
rect -536 -178 -518 -174
rect -484 -178 -466 -174
rect -804 -188 -754 -183
rect -827 -193 -819 -189
rect -867 -307 -863 -193
rect -827 -204 -823 -193
rect -839 -216 -835 -211
rect -839 -219 -831 -216
rect -867 -311 -822 -307
rect -863 -403 -858 -311
rect -825 -338 -822 -311
rect -809 -312 -806 -211
rect -796 -278 -792 -188
rect -758 -205 -739 -201
rect -730 -207 -726 -178
rect -708 -189 -702 -185
rect -678 -187 -674 -178
rect -588 -187 -546 -183
rect -678 -188 -546 -187
rect -678 -191 -584 -188
rect -730 -211 -687 -207
rect -730 -215 -726 -211
rect -678 -215 -674 -191
rect -756 -225 -752 -221
rect -704 -225 -700 -221
rect -756 -229 -748 -225
rect -704 -229 -696 -225
rect -782 -245 -774 -242
rect -757 -245 -727 -242
rect -782 -255 -778 -245
rect -757 -255 -753 -245
rect -731 -255 -727 -245
rect -705 -245 -675 -242
rect -705 -255 -701 -245
rect -679 -255 -675 -245
rect -796 -283 -779 -278
rect -769 -279 -765 -267
rect -744 -279 -740 -267
rect -692 -279 -688 -267
rect -769 -283 -754 -279
rect -744 -283 -726 -279
rect -692 -283 -674 -279
rect -769 -294 -765 -283
rect -781 -306 -777 -301
rect -781 -309 -773 -306
rect -730 -308 -726 -283
rect -709 -300 -702 -296
rect -678 -300 -674 -283
rect -663 -280 -659 -191
rect -651 -300 -647 -200
rect -617 -205 -599 -201
rect -678 -304 -643 -300
rect -730 -312 -687 -308
rect -809 -316 -739 -312
rect -730 -320 -726 -312
rect -678 -320 -674 -304
rect -756 -330 -752 -326
rect -704 -330 -700 -326
rect -756 -334 -748 -330
rect -704 -334 -696 -330
rect -617 -338 -614 -205
rect -604 -312 -600 -205
rect -588 -278 -584 -191
rect -546 -205 -531 -201
rect -522 -207 -518 -178
rect -500 -189 -494 -185
rect -470 -187 -466 -178
rect -355 -179 -351 -68
rect -341 -90 -338 -68
rect -325 -71 -321 -68
rect -335 -84 -331 -81
rect -335 -87 -321 -84
rect -312 -89 -289 -85
rect -312 -90 -308 -89
rect -341 -93 -308 -90
rect -281 -92 -277 -68
rect -269 -71 -259 -67
rect -251 -68 -243 -64
rect -253 -84 -249 -81
rect -262 -88 -249 -84
rect -301 -96 -258 -92
rect -343 -100 -309 -96
rect -348 -172 -344 -101
rect -322 -133 -319 -100
rect -301 -106 -297 -96
rect -291 -103 -267 -99
rect -291 -106 -287 -103
rect -271 -106 -267 -103
rect -311 -119 -307 -116
rect -291 -119 -287 -116
rect -311 -123 -287 -119
rect -281 -126 -277 -116
rect -313 -130 -266 -126
rect -246 -133 -243 -68
rect -239 -86 -235 -62
rect -89 -65 -49 -61
rect 45 -58 62 -53
rect -182 -71 -144 -66
rect -182 -80 -177 -71
rect -158 -80 -154 -71
rect -239 -89 -201 -86
rect -239 -91 -235 -89
rect -204 -119 -201 -89
rect -148 -80 -144 -71
rect 0 -68 34 -64
rect -167 -100 -163 -91
rect -189 -106 -179 -103
rect -167 -104 -155 -100
rect -159 -108 -144 -104
rect -136 -106 -132 -91
rect -90 -91 -38 -87
rect -90 -101 -84 -91
rect -43 -101 -38 -91
rect -204 -122 -166 -119
rect -322 -136 -243 -133
rect -237 -135 -226 -131
rect -159 -132 -155 -108
rect -136 -110 -104 -106
rect -136 -131 -132 -110
rect -107 -124 -104 -110
rect -107 -128 -85 -124
rect -56 -126 -51 -112
rect -341 -143 -287 -139
rect -335 -146 -331 -143
rect -315 -146 -311 -143
rect -307 -146 -303 -143
rect -237 -155 -233 -135
rect -56 -131 -39 -126
rect -30 -129 -26 -112
rect 0 -129 4 -68
rect 45 -84 50 -58
rect 29 -89 50 -84
rect 71 -60 75 -39
rect 97 -58 126 -54
rect 135 -56 139 -38
rect 173 -55 177 -38
rect 97 -60 101 -58
rect 71 -64 101 -60
rect 29 -92 34 -89
rect 71 -92 75 -64
rect 112 -86 116 -58
rect 135 -60 163 -56
rect 173 -59 190 -55
rect 215 -56 219 -38
rect 135 -68 139 -60
rect 149 -72 177 -68
rect 123 -80 127 -77
rect 123 -83 134 -80
rect 149 -86 153 -72
rect 112 -89 153 -86
rect 186 -88 190 -59
rect 200 -60 219 -56
rect 228 -60 240 -56
rect 215 -67 219 -60
rect 227 -79 231 -76
rect 223 -83 231 -79
rect 14 -108 19 -100
rect 45 -108 50 -100
rect 160 -92 201 -88
rect 137 -98 151 -94
rect 60 -108 65 -100
rect 14 -113 65 -108
rect -181 -145 -177 -140
rect -145 -145 -141 -139
rect -181 -149 -141 -145
rect -99 -142 -67 -138
rect -99 -161 -95 -142
rect -56 -157 -51 -131
rect -325 -172 -321 -166
rect -348 -176 -333 -172
rect -325 -176 -311 -172
rect -315 -179 -311 -176
rect -297 -179 -293 -166
rect -230 -163 -95 -161
rect -230 -164 -182 -163
rect -230 -179 -227 -164
rect -177 -164 -95 -163
rect -72 -162 -51 -157
rect -30 -133 4 -129
rect 137 -132 141 -98
rect 160 -104 164 -92
rect 172 -100 204 -95
rect 172 -104 177 -100
rect 199 -104 204 -100
rect 147 -119 152 -114
rect 172 -119 177 -114
rect 147 -123 177 -119
rect 186 -125 190 -114
rect 180 -129 190 -125
rect 236 -131 240 -60
rect 266 -129 271 -38
rect 307 -65 310 -38
rect 323 -39 326 62
rect 336 -5 340 85
rect 374 68 393 72
rect 402 66 406 95
rect 424 84 430 88
rect 454 86 458 95
rect 544 86 586 90
rect 454 85 586 86
rect 454 82 548 85
rect 402 62 445 66
rect 402 58 406 62
rect 454 58 458 82
rect 376 48 380 52
rect 428 48 432 52
rect 376 44 384 48
rect 428 44 436 48
rect 350 28 358 31
rect 375 28 405 31
rect 350 18 354 28
rect 375 18 379 28
rect 401 18 405 28
rect 427 28 457 31
rect 427 18 431 28
rect 453 18 457 28
rect 336 -10 353 -5
rect 363 -6 367 6
rect 388 -6 392 6
rect 440 -6 444 6
rect 363 -10 378 -6
rect 388 -10 406 -6
rect 440 -10 458 -6
rect 363 -21 367 -10
rect 351 -33 355 -28
rect 351 -36 359 -33
rect 402 -35 406 -10
rect 423 -27 430 -23
rect 454 -27 458 -10
rect 469 -7 473 82
rect 481 -27 485 73
rect 515 68 533 72
rect 454 -31 489 -27
rect 402 -39 445 -35
rect 323 -43 393 -39
rect 402 -47 406 -39
rect 454 -47 458 -31
rect 376 -57 380 -53
rect 428 -57 432 -53
rect 376 -61 384 -57
rect 428 -61 436 -57
rect 515 -65 518 68
rect 528 -39 532 68
rect 544 -5 548 82
rect 586 68 601 72
rect 610 66 614 95
rect 632 84 638 88
rect 662 86 666 95
rect 662 82 706 86
rect 610 62 653 66
rect 610 58 614 62
rect 662 58 666 82
rect 584 48 588 52
rect 636 48 640 52
rect 584 44 592 48
rect 636 44 644 48
rect 558 28 566 31
rect 583 28 613 31
rect 558 18 562 28
rect 583 18 587 28
rect 609 18 613 28
rect 635 28 665 31
rect 635 18 639 28
rect 661 18 665 28
rect 544 -10 561 -5
rect 571 -6 575 6
rect 596 -6 600 6
rect 648 -6 652 6
rect 571 -10 586 -6
rect 596 -10 614 -6
rect 648 -10 666 -6
rect 571 -21 575 -10
rect 559 -33 563 -28
rect 559 -36 567 -33
rect 610 -35 614 -10
rect 631 -27 638 -23
rect 662 -27 666 -10
rect 677 -7 681 82
rect 689 -27 693 73
rect 662 -31 697 -27
rect 610 -39 653 -35
rect 528 -43 601 -39
rect 610 -47 614 -39
rect 662 -47 666 -31
rect 584 -57 588 -53
rect 636 -57 640 -53
rect 584 -61 592 -57
rect 636 -61 644 -57
rect 307 -69 518 -65
rect 369 -81 399 -78
rect 369 -91 373 -81
rect 395 -91 399 -81
rect 286 -96 294 -93
rect 286 -106 290 -96
rect 421 -81 451 -78
rect 421 -91 425 -81
rect 447 -91 451 -81
rect 577 -81 607 -78
rect 577 -91 581 -81
rect 603 -91 607 -81
rect 629 -81 659 -78
rect 629 -91 633 -81
rect 655 -91 659 -81
rect 222 -132 240 -131
rect -72 -165 -67 -162
rect -30 -165 -26 -133
rect 137 -136 240 -132
rect 259 -134 289 -129
rect 299 -130 303 -118
rect 382 -115 386 -103
rect 434 -115 438 -103
rect 590 -115 594 -103
rect 642 -115 646 -103
rect 382 -119 400 -115
rect 434 -119 452 -115
rect 590 -119 608 -115
rect 642 -119 660 -115
rect 322 -129 372 -124
rect 299 -134 307 -130
rect 137 -148 140 -136
rect -355 -183 -323 -179
rect -315 -183 -305 -179
rect -297 -183 -227 -179
rect -87 -181 -82 -173
rect -56 -181 -51 -173
rect -9 -153 140 -148
rect -9 -163 -5 -153
rect -41 -181 -36 -173
rect -315 -186 -311 -183
rect -297 -186 -293 -183
rect -470 -191 -353 -187
rect -522 -211 -479 -207
rect -522 -215 -518 -211
rect -470 -215 -466 -191
rect -548 -225 -544 -221
rect -496 -225 -492 -221
rect -548 -229 -540 -225
rect -496 -229 -488 -225
rect -574 -245 -566 -242
rect -549 -245 -519 -242
rect -574 -255 -570 -245
rect -549 -255 -545 -245
rect -523 -255 -519 -245
rect -497 -245 -467 -242
rect -497 -255 -493 -245
rect -471 -255 -467 -245
rect -588 -283 -571 -278
rect -561 -279 -557 -267
rect -536 -279 -532 -267
rect -484 -279 -480 -267
rect -561 -283 -546 -279
rect -536 -283 -518 -279
rect -484 -283 -466 -279
rect -561 -294 -557 -283
rect -573 -306 -569 -301
rect -573 -309 -565 -306
rect -522 -308 -518 -283
rect -501 -300 -494 -296
rect -470 -300 -466 -283
rect -455 -280 -451 -191
rect -443 -300 -439 -200
rect -356 -242 -353 -191
rect -154 -190 -116 -185
rect -87 -186 -36 -181
rect -335 -199 -331 -196
rect -307 -199 -303 -196
rect -154 -199 -149 -190
rect -130 -199 -126 -190
rect -341 -203 -282 -199
rect -341 -213 -243 -209
rect -120 -199 -116 -190
rect -335 -216 -331 -213
rect -311 -216 -307 -213
rect -271 -216 -267 -213
rect -253 -216 -249 -213
rect -139 -219 -135 -210
rect -190 -224 -151 -221
rect -139 -223 -127 -219
rect -131 -227 -116 -223
rect -108 -225 -104 -210
rect -71 -204 -33 -199
rect -71 -213 -66 -204
rect -47 -213 -43 -204
rect -37 -213 -33 -204
rect 12 -212 50 -207
rect -325 -242 -321 -236
rect -291 -242 -287 -236
rect -359 -246 -333 -242
rect -325 -246 -299 -242
rect -291 -246 -277 -242
rect -263 -245 -259 -236
rect -211 -242 -138 -238
rect -470 -304 -435 -300
rect -522 -312 -479 -308
rect -604 -316 -531 -312
rect -522 -320 -518 -312
rect -470 -320 -466 -304
rect -548 -330 -544 -326
rect -496 -330 -492 -326
rect -548 -334 -540 -330
rect -496 -334 -488 -330
rect -825 -342 -614 -338
rect -766 -355 -736 -352
rect -766 -365 -762 -355
rect -740 -365 -736 -355
rect -849 -370 -841 -367
rect -849 -380 -845 -370
rect -714 -355 -684 -352
rect -714 -365 -710 -355
rect -688 -365 -684 -355
rect -558 -355 -528 -352
rect -558 -365 -554 -355
rect -532 -365 -528 -355
rect -506 -355 -476 -352
rect -506 -365 -502 -355
rect -480 -365 -476 -355
rect -876 -408 -846 -403
rect -836 -404 -832 -392
rect -753 -389 -749 -377
rect -701 -389 -697 -377
rect -545 -389 -541 -377
rect -493 -389 -489 -377
rect -753 -393 -735 -389
rect -701 -393 -683 -389
rect -545 -393 -527 -389
rect -493 -393 -475 -389
rect -813 -403 -763 -398
rect -836 -408 -828 -404
rect -876 -522 -872 -408
rect -836 -419 -832 -408
rect -848 -431 -844 -426
rect -848 -434 -840 -431
rect -876 -526 -831 -522
rect -834 -553 -831 -526
rect -818 -527 -815 -426
rect -805 -493 -801 -403
rect -767 -420 -748 -416
rect -739 -422 -735 -393
rect -717 -404 -711 -400
rect -687 -402 -683 -393
rect -597 -402 -555 -398
rect -687 -403 -555 -402
rect -687 -406 -593 -403
rect -739 -426 -696 -422
rect -739 -430 -735 -426
rect -687 -430 -683 -406
rect -765 -440 -761 -436
rect -713 -440 -709 -436
rect -765 -444 -757 -440
rect -713 -444 -705 -440
rect -791 -460 -783 -457
rect -766 -460 -736 -457
rect -791 -470 -787 -460
rect -766 -470 -762 -460
rect -740 -470 -736 -460
rect -714 -460 -684 -457
rect -714 -470 -710 -460
rect -688 -470 -684 -460
rect -805 -498 -788 -493
rect -778 -494 -774 -482
rect -753 -494 -749 -482
rect -701 -494 -697 -482
rect -778 -498 -763 -494
rect -753 -498 -735 -494
rect -701 -498 -683 -494
rect -778 -509 -774 -498
rect -790 -521 -786 -516
rect -790 -524 -782 -521
rect -739 -523 -735 -498
rect -718 -515 -711 -511
rect -687 -515 -683 -498
rect -672 -495 -668 -406
rect -660 -515 -656 -415
rect -626 -420 -608 -416
rect -687 -519 -652 -515
rect -739 -527 -696 -523
rect -818 -531 -748 -527
rect -739 -535 -735 -527
rect -687 -535 -683 -519
rect -765 -545 -761 -541
rect -713 -545 -709 -541
rect -765 -549 -757 -545
rect -713 -549 -705 -545
rect -626 -553 -623 -420
rect -613 -527 -609 -420
rect -597 -493 -593 -406
rect -555 -420 -540 -416
rect -531 -422 -527 -393
rect -509 -404 -503 -400
rect -479 -402 -475 -393
rect -406 -402 -402 -275
rect -355 -357 -351 -246
rect -341 -268 -338 -246
rect -325 -249 -321 -246
rect -335 -262 -331 -259
rect -335 -265 -321 -262
rect -312 -267 -289 -263
rect -312 -268 -308 -267
rect -341 -271 -308 -268
rect -281 -270 -277 -246
rect -269 -249 -259 -245
rect -251 -246 -243 -242
rect -253 -262 -249 -259
rect -262 -266 -249 -262
rect -301 -274 -258 -270
rect -343 -278 -309 -274
rect -348 -350 -344 -279
rect -322 -311 -319 -278
rect -301 -284 -297 -274
rect -291 -281 -267 -277
rect -291 -284 -287 -281
rect -271 -284 -267 -281
rect -311 -297 -307 -294
rect -291 -297 -287 -294
rect -311 -301 -287 -297
rect -281 -304 -277 -294
rect -313 -308 -266 -304
rect -246 -311 -243 -246
rect -131 -251 -127 -227
rect -108 -229 -86 -225
rect -108 -250 -104 -229
rect -89 -235 -86 -229
rect -56 -233 -52 -224
rect -89 -238 -68 -235
rect -56 -237 -44 -233
rect -48 -241 -33 -237
rect -25 -239 -21 -224
rect 12 -221 17 -212
rect 36 -221 40 -212
rect 46 -221 50 -212
rect -88 -255 -55 -252
rect -153 -264 -149 -259
rect -117 -264 -113 -258
rect -153 -268 -113 -264
rect -48 -265 -44 -241
rect -25 -243 -10 -239
rect 27 -241 31 -232
rect -25 -264 -21 -243
rect -13 -247 15 -243
rect 27 -245 39 -241
rect 35 -249 50 -245
rect 58 -247 62 -232
rect -233 -275 -229 -270
rect -232 -292 -229 -275
rect 3 -264 28 -260
rect -70 -278 -66 -273
rect -34 -278 -30 -272
rect -70 -282 -30 -278
rect 3 -292 6 -264
rect 35 -273 39 -249
rect 58 -251 73 -247
rect 259 -248 263 -134
rect 299 -145 303 -134
rect 287 -157 291 -152
rect 287 -160 295 -157
rect 58 -272 62 -251
rect 13 -286 17 -281
rect 49 -286 53 -280
rect 13 -290 53 -286
rect 69 -286 73 -251
rect 91 -254 143 -250
rect 259 -252 304 -248
rect 91 -264 97 -254
rect 138 -264 143 -254
rect 301 -259 304 -252
rect 317 -253 320 -152
rect 330 -219 334 -129
rect 368 -146 387 -142
rect 396 -148 400 -119
rect 418 -130 424 -126
rect 448 -128 452 -119
rect 538 -128 580 -124
rect 448 -129 580 -128
rect 448 -132 542 -129
rect 396 -152 439 -148
rect 396 -156 400 -152
rect 448 -156 452 -132
rect 370 -166 374 -162
rect 422 -166 426 -162
rect 370 -170 378 -166
rect 422 -170 430 -166
rect 344 -186 352 -183
rect 369 -186 399 -183
rect 344 -196 348 -186
rect 369 -196 373 -186
rect 395 -196 399 -186
rect 421 -186 451 -183
rect 421 -196 425 -186
rect 447 -196 451 -186
rect 330 -224 347 -219
rect 357 -220 361 -208
rect 382 -220 386 -208
rect 434 -220 438 -208
rect 357 -224 372 -220
rect 382 -224 400 -220
rect 434 -224 452 -220
rect 357 -235 361 -224
rect 345 -247 349 -242
rect 345 -250 353 -247
rect 396 -249 400 -224
rect 417 -241 424 -237
rect 448 -241 452 -224
rect 463 -221 467 -132
rect 475 -241 479 -141
rect 509 -146 527 -142
rect 448 -245 483 -241
rect 396 -253 439 -249
rect 317 -257 387 -253
rect 187 -260 304 -259
rect 69 -291 96 -286
rect 125 -289 130 -275
rect -232 -294 6 -292
rect -232 -296 -75 -294
rect -70 -296 6 -294
rect 125 -294 142 -289
rect -322 -314 -243 -311
rect -139 -306 -101 -301
rect -139 -315 -134 -306
rect -115 -315 -111 -306
rect -341 -321 -287 -317
rect -335 -324 -331 -321
rect -315 -324 -311 -321
rect -307 -324 -303 -321
rect -105 -315 -101 -306
rect 54 -305 114 -301
rect -325 -350 -321 -344
rect -348 -354 -333 -350
rect -325 -354 -311 -350
rect -315 -357 -311 -354
rect -297 -357 -293 -344
rect -124 -335 -120 -326
rect -228 -343 -223 -339
rect -164 -341 -136 -338
rect -124 -339 -112 -335
rect -164 -343 -161 -341
rect -228 -346 -161 -343
rect -116 -343 -101 -339
rect -93 -341 -89 -326
rect -56 -320 -18 -315
rect -56 -329 -51 -320
rect -32 -329 -28 -320
rect -22 -329 -18 -320
rect -355 -361 -323 -357
rect -315 -361 -305 -357
rect -297 -361 -228 -357
rect -196 -358 -123 -354
rect -315 -364 -311 -361
rect -297 -364 -293 -361
rect -335 -377 -331 -374
rect -307 -377 -303 -374
rect -341 -381 -282 -377
rect -479 -406 -402 -402
rect -531 -426 -488 -422
rect -531 -430 -527 -426
rect -479 -430 -475 -406
rect -557 -440 -553 -436
rect -505 -440 -501 -436
rect -557 -444 -549 -440
rect -505 -444 -497 -440
rect -583 -460 -575 -457
rect -558 -460 -528 -457
rect -583 -470 -579 -460
rect -558 -470 -554 -460
rect -532 -470 -528 -460
rect -506 -460 -476 -457
rect -506 -470 -502 -460
rect -480 -470 -476 -460
rect -597 -498 -580 -493
rect -570 -494 -566 -482
rect -545 -494 -541 -482
rect -493 -494 -489 -482
rect -570 -498 -555 -494
rect -545 -498 -527 -494
rect -493 -498 -475 -494
rect -570 -509 -566 -498
rect -582 -521 -578 -516
rect -582 -524 -574 -521
rect -531 -523 -527 -498
rect -510 -515 -503 -511
rect -479 -515 -475 -498
rect -464 -495 -460 -406
rect -452 -515 -448 -415
rect -232 -492 -228 -361
rect -116 -367 -112 -343
rect -93 -345 -71 -341
rect -93 -366 -89 -345
rect -74 -351 -71 -345
rect -41 -349 -37 -340
rect -10 -348 -6 -340
rect 54 -348 58 -305
rect 125 -320 130 -294
rect 109 -325 130 -320
rect 151 -321 155 -275
rect 183 -265 304 -260
rect 396 -261 400 -253
rect 448 -261 452 -245
rect 151 -325 165 -321
rect 109 -328 114 -325
rect 151 -328 155 -325
rect -74 -354 -53 -351
rect -41 -353 -29 -349
rect -10 -352 58 -348
rect 94 -344 99 -336
rect 125 -344 130 -336
rect 140 -344 145 -336
rect 94 -349 145 -344
rect -33 -357 -18 -353
rect -65 -372 -40 -369
rect -138 -380 -134 -375
rect -102 -380 -98 -374
rect -138 -384 -98 -380
rect -33 -381 -29 -357
rect -10 -380 -6 -352
rect 161 -359 165 -325
rect 183 -353 188 -265
rect 301 -279 304 -265
rect 370 -271 374 -267
rect 422 -271 426 -267
rect 370 -275 378 -271
rect 422 -275 430 -271
rect 509 -279 512 -146
rect 522 -253 526 -146
rect 538 -219 542 -132
rect 580 -146 595 -142
rect 604 -148 608 -119
rect 626 -130 632 -126
rect 656 -128 660 -119
rect 656 -132 693 -128
rect 604 -152 647 -148
rect 604 -156 608 -152
rect 656 -156 660 -132
rect 578 -166 582 -162
rect 630 -166 634 -162
rect 578 -170 586 -166
rect 630 -170 638 -166
rect 552 -186 560 -183
rect 577 -186 607 -183
rect 552 -196 556 -186
rect 577 -196 581 -186
rect 603 -196 607 -186
rect 629 -186 659 -183
rect 629 -196 633 -186
rect 655 -196 659 -186
rect 538 -224 555 -219
rect 565 -220 569 -208
rect 590 -220 594 -208
rect 642 -220 646 -208
rect 565 -224 580 -220
rect 590 -224 608 -220
rect 642 -224 660 -220
rect 565 -235 569 -224
rect 553 -247 557 -242
rect 553 -250 561 -247
rect 604 -249 608 -224
rect 625 -241 632 -237
rect 656 -241 660 -224
rect 671 -221 675 -132
rect 683 -241 687 -141
rect 656 -245 691 -241
rect 604 -253 647 -249
rect 522 -257 595 -253
rect 604 -261 608 -253
rect 656 -261 660 -245
rect 578 -271 582 -267
rect 630 -271 634 -267
rect 578 -275 586 -271
rect 630 -275 638 -271
rect 301 -283 512 -279
rect 282 -305 312 -302
rect 282 -315 286 -305
rect 308 -315 312 -305
rect 199 -320 207 -317
rect 199 -330 203 -320
rect 334 -305 364 -302
rect 334 -315 338 -305
rect 360 -315 364 -305
rect 490 -305 520 -302
rect 490 -315 494 -305
rect 516 -315 520 -305
rect 542 -305 572 -302
rect 542 -315 546 -305
rect 568 -315 572 -305
rect 37 -363 165 -359
rect 172 -358 202 -353
rect 212 -354 216 -342
rect 295 -339 299 -327
rect 347 -339 351 -327
rect 503 -339 507 -327
rect 555 -339 559 -327
rect 295 -343 313 -339
rect 347 -343 365 -339
rect 503 -343 521 -339
rect 555 -343 573 -339
rect 235 -353 285 -348
rect 212 -358 220 -354
rect -55 -394 -51 -389
rect -19 -394 -15 -388
rect -141 -400 -103 -395
rect -55 -398 -15 -394
rect -141 -409 -136 -400
rect -117 -409 -113 -400
rect -107 -409 -103 -400
rect 37 -404 42 -363
rect 55 -371 107 -367
rect 55 -381 61 -371
rect 102 -381 107 -371
rect 37 -408 60 -404
rect 89 -406 94 -392
rect -126 -429 -122 -420
rect -173 -435 -138 -431
rect -126 -433 -114 -429
rect -118 -437 -103 -433
rect -95 -435 -91 -420
rect -46 -414 6 -410
rect -46 -424 -40 -414
rect 1 -424 6 -414
rect 89 -411 106 -406
rect 45 -422 78 -418
rect -212 -451 -125 -448
rect -118 -461 -114 -437
rect -95 -439 -67 -435
rect -95 -460 -91 -439
rect -71 -447 -67 -439
rect -71 -451 -41 -447
rect -12 -449 -7 -435
rect -12 -454 5 -449
rect -60 -465 -23 -460
rect -140 -474 -136 -469
rect -104 -474 -100 -468
rect -140 -478 -100 -474
rect -60 -492 -56 -465
rect -12 -480 -7 -454
rect -28 -485 -7 -480
rect 14 -459 18 -435
rect 45 -459 49 -422
rect 89 -437 94 -411
rect 73 -442 94 -437
rect 115 -419 119 -392
rect 115 -424 130 -419
rect 73 -445 78 -442
rect 115 -445 119 -424
rect 14 -464 49 -459
rect 58 -461 63 -453
rect 89 -461 94 -453
rect 104 -461 109 -453
rect -28 -488 -23 -485
rect 14 -488 18 -464
rect 58 -466 109 -461
rect 172 -472 176 -358
rect 212 -369 216 -358
rect 200 -381 204 -376
rect 200 -384 208 -381
rect 172 -476 217 -472
rect -232 -497 -56 -492
rect -43 -504 -38 -496
rect -12 -504 -7 -496
rect 3 -504 8 -496
rect -43 -509 8 -504
rect 214 -503 217 -476
rect 230 -477 233 -376
rect 243 -443 247 -353
rect 281 -370 300 -366
rect 309 -372 313 -343
rect 331 -354 337 -350
rect 361 -352 365 -343
rect 451 -352 493 -348
rect 361 -353 493 -352
rect 361 -356 455 -353
rect 309 -376 352 -372
rect 309 -380 313 -376
rect 361 -380 365 -356
rect 283 -390 287 -386
rect 335 -390 339 -386
rect 283 -394 291 -390
rect 335 -394 343 -390
rect 257 -410 265 -407
rect 282 -410 312 -407
rect 257 -420 261 -410
rect 282 -420 286 -410
rect 308 -420 312 -410
rect 334 -410 364 -407
rect 334 -420 338 -410
rect 360 -420 364 -410
rect 243 -448 260 -443
rect 270 -444 274 -432
rect 295 -444 299 -432
rect 347 -444 351 -432
rect 270 -448 285 -444
rect 295 -448 313 -444
rect 347 -448 365 -444
rect 270 -459 274 -448
rect 258 -471 262 -466
rect 258 -474 266 -471
rect 309 -473 313 -448
rect 330 -465 337 -461
rect 361 -465 365 -448
rect 376 -445 380 -356
rect 388 -465 392 -365
rect 422 -370 440 -366
rect 361 -469 396 -465
rect 309 -477 352 -473
rect 230 -481 300 -477
rect 309 -485 313 -477
rect 361 -485 365 -469
rect 283 -495 287 -491
rect 335 -495 339 -491
rect 283 -499 291 -495
rect 335 -499 343 -495
rect 422 -503 425 -370
rect 435 -477 439 -370
rect 451 -443 455 -356
rect 493 -370 508 -366
rect 517 -372 521 -343
rect 539 -354 545 -350
rect 569 -352 573 -343
rect 569 -356 605 -352
rect 517 -376 560 -372
rect 517 -380 521 -376
rect 569 -380 573 -356
rect 491 -390 495 -386
rect 543 -390 547 -386
rect 491 -394 499 -390
rect 543 -394 551 -390
rect 465 -410 473 -407
rect 490 -410 520 -407
rect 465 -420 469 -410
rect 490 -420 494 -410
rect 516 -420 520 -410
rect 542 -410 572 -407
rect 542 -420 546 -410
rect 568 -420 572 -410
rect 451 -448 468 -443
rect 478 -444 482 -432
rect 503 -444 507 -432
rect 555 -444 559 -432
rect 478 -448 493 -444
rect 503 -448 521 -444
rect 555 -448 573 -444
rect 478 -459 482 -448
rect 466 -471 470 -466
rect 466 -474 474 -471
rect 517 -473 521 -448
rect 538 -465 545 -461
rect 569 -465 573 -448
rect 584 -445 588 -356
rect 596 -465 600 -365
rect 569 -469 604 -465
rect 517 -477 560 -473
rect 435 -481 508 -477
rect 517 -485 521 -477
rect 569 -485 573 -469
rect 491 -495 495 -491
rect 543 -495 547 -491
rect 491 -499 499 -495
rect 543 -499 551 -495
rect 214 -507 425 -503
rect -479 -519 -444 -515
rect -531 -527 -488 -523
rect -613 -531 -540 -527
rect -531 -535 -527 -527
rect -479 -535 -475 -519
rect -557 -545 -553 -541
rect -505 -545 -501 -541
rect -557 -549 -549 -545
rect -505 -549 -497 -545
rect -834 -557 -623 -553
<< m2contact >>
rect -813 728 -808 733
rect -831 720 -826 725
rect -825 672 -820 677
rect -921 623 -915 628
rect -809 622 -804 627
rect -905 572 -900 577
rect -825 508 -820 513
rect -568 719 -563 724
rect -586 711 -581 716
rect -580 663 -575 668
rect -676 614 -670 619
rect -564 613 -559 618
rect -660 563 -655 568
rect -825 460 -820 465
rect -580 499 -575 504
rect -307 743 -302 748
rect -325 735 -320 740
rect -319 687 -314 692
rect -415 638 -409 643
rect -303 637 -298 642
rect -399 587 -394 592
rect -921 415 -915 420
rect -580 451 -575 456
rect -319 523 -314 528
rect -319 475 -314 480
rect -182 512 -177 517
rect -235 504 -230 509
rect -809 414 -804 419
rect -676 406 -670 411
rect -564 405 -559 410
rect -415 430 -409 435
rect -303 429 -298 434
rect -174 494 -169 499
rect -399 379 -394 384
rect -905 364 -900 369
rect -931 281 -926 286
rect -949 273 -944 278
rect -943 225 -938 230
rect -660 355 -655 360
rect -126 500 -121 505
rect -76 516 -71 521
rect -163 460 -158 465
rect -77 404 -72 410
rect -26 420 -21 425
rect 38 500 43 505
rect 86 500 91 505
rect 132 516 137 521
rect 131 404 136 410
rect 182 420 187 425
rect -373 342 -368 347
rect -804 252 -799 257
rect -1039 176 -1033 181
rect -927 175 -922 180
rect -1023 125 -1018 130
rect -943 61 -938 66
rect -796 234 -791 239
rect -943 13 -938 18
rect -748 240 -743 245
rect -698 256 -693 261
rect -699 144 -694 150
rect -648 160 -643 165
rect -584 240 -579 245
rect -536 240 -531 245
rect -490 256 -485 261
rect -491 144 -486 150
rect -440 160 -435 165
rect -395 110 -390 115
rect 92 307 97 312
rect -348 255 -343 260
rect -258 259 -252 265
rect -219 268 -214 274
rect -98 235 -93 240
rect 100 289 105 294
rect -203 132 -198 137
rect 110 245 115 251
rect 148 295 153 300
rect 198 311 203 316
rect 197 199 202 205
rect 248 215 253 220
rect 312 295 317 300
rect 360 295 365 300
rect 406 311 411 316
rect 405 199 410 205
rect 456 215 461 220
rect -224 120 -219 126
rect -817 38 -812 43
rect -1039 -32 -1033 -27
rect -927 -33 -922 -28
rect -1023 -83 -1018 -78
rect -809 20 -804 25
rect -761 26 -756 31
rect -711 42 -706 47
rect -712 -70 -707 -64
rect -661 -54 -656 -49
rect -597 26 -592 31
rect -549 26 -544 31
rect -503 42 -498 47
rect -504 -70 -499 -64
rect -453 -54 -448 -49
rect -348 77 -343 82
rect -258 81 -252 87
rect -236 82 -231 87
rect 141 69 146 74
rect -98 40 -93 46
rect -203 32 -198 39
rect 313 80 318 85
rect -234 -36 -228 -30
rect -178 -24 -173 -19
rect -103 -36 -98 -31
rect -215 -51 -210 -46
rect 321 62 326 67
rect -420 -115 -415 -110
rect -819 -193 -814 -188
rect -811 -211 -806 -206
rect -763 -205 -758 -200
rect -713 -189 -708 -184
rect -714 -301 -709 -295
rect -663 -285 -658 -280
rect -599 -205 -594 -200
rect -551 -205 -546 -200
rect -505 -189 -500 -184
rect -348 -101 -343 -96
rect -258 -97 -252 -91
rect -240 -96 -235 -91
rect -195 -106 -189 -101
rect -226 -135 -221 -130
rect 201 -92 206 -87
rect -238 -160 -233 -155
rect -182 -168 -177 -163
rect 331 45 336 51
rect 369 68 374 73
rect 419 84 424 89
rect 418 -28 423 -22
rect 469 -12 474 -7
rect 533 68 538 73
rect 581 68 586 73
rect 627 84 632 89
rect 626 -28 631 -22
rect 677 -12 682 -7
rect 307 -134 312 -129
rect -9 -169 -4 -163
rect -506 -301 -501 -295
rect -455 -285 -450 -280
rect -195 -224 -190 -219
rect -216 -242 -211 -237
rect -828 -408 -823 -403
rect -820 -426 -815 -421
rect -772 -420 -767 -415
rect -722 -404 -717 -399
rect -723 -516 -718 -510
rect -672 -500 -667 -495
rect -608 -420 -603 -415
rect -560 -420 -555 -415
rect -514 -404 -509 -399
rect -402 -279 -397 -274
rect -348 -279 -343 -274
rect -258 -275 -252 -269
rect -93 -255 -88 -250
rect -238 -275 -233 -269
rect -9 -292 -4 -287
rect 315 -152 320 -147
rect 324 -182 330 -175
rect 363 -146 368 -141
rect 413 -130 418 -125
rect 412 -242 417 -236
rect 463 -226 468 -221
rect 527 -146 532 -141
rect -217 -301 -212 -296
rect -75 -299 -70 -294
rect -228 -339 -223 -334
rect -201 -359 -196 -354
rect -515 -516 -510 -510
rect -464 -500 -459 -495
rect -70 -372 -65 -367
rect 575 -146 580 -141
rect 621 -130 626 -125
rect 620 -242 625 -236
rect 671 -226 676 -221
rect 220 -358 225 -353
rect -218 -451 -212 -445
rect 130 -425 136 -418
rect 228 -376 233 -371
rect 238 -424 243 -419
rect 276 -370 281 -365
rect 326 -354 331 -349
rect 325 -466 330 -460
rect 376 -450 381 -445
rect 440 -370 445 -365
rect 488 -370 493 -365
rect 534 -354 539 -349
rect 533 -466 538 -460
rect 584 -450 589 -445
<< pdm12contact >>
rect -820 560 -815 565
rect -575 551 -570 556
rect -314 575 -309 580
rect -820 352 -815 357
rect -314 367 -309 372
rect -14 505 -9 510
rect 194 505 199 510
rect -575 343 -570 348
rect -938 113 -933 118
rect -636 245 -631 250
rect -428 245 -423 250
rect 260 300 265 305
rect 468 300 473 305
rect -938 -95 -933 -90
rect -649 31 -644 36
rect -441 31 -436 36
rect -651 -200 -646 -195
rect 481 73 486 78
rect 689 73 694 78
rect -443 -200 -438 -195
rect -660 -415 -655 -410
rect 475 -141 480 -136
rect -452 -415 -447 -410
rect 683 -141 688 -136
rect -178 -435 -173 -430
rect 388 -365 393 -360
rect 596 -365 601 -360
<< metal2 >>
rect -325 744 -307 747
rect -325 740 -321 744
rect -831 729 -813 732
rect -831 725 -827 729
rect -586 720 -568 723
rect -831 681 -827 720
rect -586 716 -582 720
rect -831 677 -821 681
rect -586 672 -582 711
rect -325 696 -321 735
rect -325 692 -315 696
rect -586 668 -576 672
rect -409 638 -399 642
rect -915 623 -905 627
rect -909 572 -905 623
rect -815 622 -809 626
rect -815 561 -811 622
rect -670 614 -660 618
rect -664 563 -660 614
rect -570 613 -564 617
rect -570 552 -566 613
rect -403 587 -399 638
rect -309 637 -303 641
rect -309 576 -305 637
rect -319 508 -315 523
rect -75 514 -71 516
rect 133 514 137 516
rect -825 465 -821 508
rect -319 504 -235 508
rect -580 456 -576 499
rect -319 480 -315 504
rect -181 498 -178 512
rect -75 510 -10 514
rect 133 510 198 514
rect -181 494 -174 498
rect -130 498 -126 504
rect 43 500 86 504
rect -169 494 -126 498
rect -202 460 -163 464
rect -409 430 -399 434
rect -915 415 -905 419
rect -909 364 -905 415
rect -815 414 -809 418
rect -815 353 -811 414
rect -670 406 -660 410
rect -664 355 -660 406
rect -570 405 -564 409
rect -570 344 -566 405
rect -403 379 -399 430
rect -309 429 -303 433
rect -309 368 -305 429
rect -202 387 -198 460
rect -76 416 -21 420
rect 132 416 187 420
rect -76 410 -72 416
rect 132 410 136 416
rect -240 382 -198 387
rect -949 282 -931 285
rect -949 278 -945 282
rect -949 234 -945 273
rect -373 260 -370 342
rect -373 256 -348 260
rect -697 254 -693 256
rect -489 254 -485 256
rect -240 264 -235 382
rect 199 309 203 311
rect 407 309 411 311
rect 93 293 96 307
rect 199 305 264 309
rect 407 305 472 309
rect 93 289 100 293
rect 144 293 148 299
rect 317 295 360 299
rect 105 289 148 293
rect -252 260 -235 264
rect -803 238 -800 252
rect -697 250 -632 254
rect -489 250 -424 254
rect -803 234 -796 238
rect -752 238 -748 244
rect -579 240 -536 244
rect -791 234 -748 238
rect -949 230 -939 234
rect -1033 176 -1023 180
rect -1027 125 -1023 176
rect -933 175 -927 179
rect -933 114 -929 175
rect -698 156 -643 160
rect -490 156 -435 160
rect -698 150 -694 156
rect -490 150 -486 156
rect -224 126 -219 273
rect -54 250 -50 251
rect -54 245 110 250
rect -54 239 -50 245
rect -93 235 -50 239
rect 198 211 253 215
rect 406 211 461 215
rect 198 205 202 211
rect 406 205 410 211
rect -394 82 -390 110
rect -394 78 -348 82
rect -252 82 -236 86
rect -943 18 -939 61
rect -710 40 -706 42
rect -502 40 -498 42
rect -816 24 -813 38
rect -710 36 -645 40
rect -502 36 -437 40
rect -816 20 -809 24
rect -765 24 -761 30
rect -592 26 -549 30
rect -804 20 -761 24
rect -241 -20 -237 82
rect -203 39 -198 132
rect 185 73 189 85
rect 420 82 424 84
rect 628 82 632 84
rect 146 69 189 73
rect 185 50 189 69
rect 314 66 317 80
rect 420 78 485 82
rect 628 78 693 82
rect 314 62 321 66
rect 365 66 369 72
rect 538 68 581 72
rect 326 62 369 66
rect 185 46 331 50
rect -241 -23 -178 -20
rect -1033 -32 -1023 -28
rect -1027 -83 -1023 -32
rect -933 -33 -927 -29
rect -933 -94 -929 -33
rect -233 -39 -228 -36
rect -233 -42 -191 -39
rect -711 -58 -656 -54
rect -503 -58 -448 -54
rect -711 -64 -707 -58
rect -503 -64 -499 -58
rect -420 -100 -348 -96
rect -420 -110 -416 -100
rect -252 -96 -240 -92
rect -248 -147 -244 -96
rect -226 -130 -222 -42
rect -214 -133 -211 -51
rect -194 -101 -191 -42
rect -186 -54 -183 -23
rect -102 -31 -98 46
rect 419 -16 474 -12
rect 627 -16 682 -12
rect 419 -22 423 -16
rect 627 -22 631 -16
rect -186 -57 -104 -54
rect -214 -136 -192 -133
rect -248 -151 -212 -147
rect -712 -191 -708 -189
rect -504 -191 -500 -189
rect -818 -207 -815 -193
rect -712 -195 -647 -191
rect -504 -195 -439 -191
rect -818 -211 -811 -207
rect -767 -207 -763 -201
rect -594 -205 -551 -201
rect -806 -211 -763 -207
rect -238 -219 -234 -160
rect -238 -223 -224 -219
rect -397 -278 -348 -274
rect -252 -274 -238 -270
rect -713 -289 -658 -285
rect -505 -289 -450 -285
rect -713 -295 -709 -289
rect -505 -295 -501 -289
rect -228 -334 -224 -223
rect -216 -229 -212 -151
rect -195 -219 -192 -136
rect -216 -233 -197 -229
rect -216 -237 -212 -233
rect -721 -406 -717 -404
rect -513 -406 -509 -404
rect -827 -422 -824 -408
rect -721 -410 -656 -406
rect -513 -410 -448 -406
rect -827 -426 -820 -422
rect -776 -422 -772 -416
rect -603 -420 -560 -416
rect -815 -426 -772 -422
rect -217 -445 -213 -301
rect -201 -354 -197 -233
rect -182 -435 -178 -168
rect -107 -184 -104 -57
rect 245 -88 249 -76
rect 206 -92 249 -88
rect -107 -187 -90 -184
rect -93 -250 -90 -187
rect -9 -287 -5 -169
rect 244 -176 249 -92
rect 414 -132 418 -130
rect 622 -132 626 -130
rect 308 -148 311 -134
rect 414 -136 479 -132
rect 622 -136 687 -132
rect 308 -152 315 -148
rect 359 -148 363 -142
rect 532 -146 575 -142
rect 320 -152 363 -148
rect 244 -181 324 -176
rect 413 -230 468 -226
rect 621 -230 676 -226
rect 413 -236 417 -230
rect 621 -236 625 -230
rect -74 -372 -70 -299
rect 327 -356 331 -354
rect 535 -356 539 -354
rect 221 -372 224 -358
rect 327 -360 392 -356
rect 535 -360 600 -356
rect 221 -376 228 -372
rect 272 -372 276 -366
rect 445 -370 488 -366
rect 233 -376 276 -372
rect 136 -424 238 -419
rect 326 -454 381 -450
rect 534 -454 589 -450
rect 326 -460 330 -454
rect 534 -460 538 -454
rect -722 -504 -667 -500
rect -514 -504 -459 -500
rect -722 -510 -718 -504
rect -514 -510 -510 -504
<< labels >>
rlabel metal1 -292 -308 -287 -304 1 gnd
rlabel metal1 -292 -130 -287 -126 1 gnd
rlabel metal1 -292 48 -287 52 1 gnd
rlabel metal1 -292 226 -287 230 1 gnd
rlabel metal1 -330 -265 -327 -262 1 gnd
rlabel metal1 -330 -87 -327 -84 1 gnd
rlabel metal1 -330 91 -327 94 1 gnd
rlabel metal1 -259 -265 -256 -262 1 gnd
rlabel metal1 -259 -87 -256 -84 1 gnd
rlabel metal1 -259 91 -256 94 1 gnd
rlabel metal1 -259 269 -256 272 1 gnd
rlabel metal1 -317 -213 -313 -209 4 vdd
rlabel metal1 -317 -35 -313 -31 4 vdd
rlabel metal1 -317 143 -313 147 4 vdd
rlabel metal1 -317 321 -313 325 4 vdd
rlabel metal1 -341 -321 -337 -317 4 vdd
rlabel metal1 -341 -143 -337 -139 4 vdd
rlabel metal1 -341 35 -337 39 4 vdd
rlabel metal1 -341 -381 -337 -377 2 gnd
rlabel metal1 -341 -203 -337 -199 2 gnd
rlabel metal1 -341 -25 -337 -21 2 gnd
rlabel metal1 -341 213 -337 217 4 vdd
rlabel metal1 -341 153 -337 157 2 gnd
rlabel metal1 -330 269 -326 272 1 gnd
rlabel metal1 -359 288 -355 292 3 a0
rlabel metal2 -362 256 -356 260 3 b0
rlabel metal1 -266 260 -262 264 1 p0
rlabel metal1 -284 173 -280 177 1 g0
rlabel metal1 -359 110 -356 114 3 a1
rlabel metal2 -359 78 -356 82 3 b1
rlabel metal2 -251 82 -247 86 1 p1
rlabel metal1 -282 -5 -276 -1 1 g1
rlabel metal2 -252 -96 -248 -92 1 p2
rlabel metal1 -359 -68 -356 -64 3 a2
rlabel metal2 -359 -100 -356 -96 3 b2
rlabel metal1 -359 -246 -356 -242 3 a3
rlabel metal1 -288 -183 -284 -179 1 g2
rlabel metal2 -359 -278 -356 -274 3 b3
rlabel metal2 -250 -274 -246 -270 1 p3
rlabel metal1 -287 -361 -283 -357 1 g3
rlabel metal1 -120 169 -114 174 5 vdd
rlabel metal1 -119 91 -114 95 1 gnd
rlabel metal1 -31 74 -25 79 1 gnd
rlabel metal1 -28 169 -17 173 5 vdd
rlabel metal1 16 121 20 126 1 c2
rlabel metal1 -61 -65 -56 -61 1 gnd
rlabel metal1 -62 13 -56 18 5 vdd
rlabel metal1 -144 -51 -139 -47 1 gnd
rlabel metal1 -145 27 -139 32 5 vdd
rlabel metal1 -154 -71 -148 -66 5 vdd
rlabel metal1 -153 -149 -148 -145 1 gnd
rlabel metal1 -70 -91 -59 -87 5 vdd
rlabel metal1 -73 -186 -67 -181 1 gnd
rlabel metal1 31 -18 42 -14 5 vdd
rlabel metal1 28 -113 34 -108 1 gnd
rlabel metal1 73 -64 78 -60 1 c3
rlabel metal1 -126 -190 -120 -185 5 vdd
rlabel metal1 -125 -268 -120 -264 1 gnd
rlabel metal1 -43 -204 -37 -199 5 vdd
rlabel metal1 -42 -282 -37 -278 1 gnd
rlabel metal1 40 -212 46 -207 5 vdd
rlabel metal1 41 -290 46 -286 1 gnd
rlabel metal1 -27 -398 -22 -394 1 gnd
rlabel metal1 -28 -320 -22 -315 5 vdd
rlabel metal1 -110 -384 -105 -380 1 gnd
rlabel metal1 -111 -306 -105 -301 5 vdd
rlabel metal1 -112 -478 -107 -474 1 gnd
rlabel metal1 -113 -400 -107 -395 5 vdd
rlabel metal1 111 -254 122 -250 5 vdd
rlabel metal1 108 -349 114 -344 1 gnd
rlabel metal1 75 -371 86 -367 5 vdd
rlabel metal1 72 -466 78 -461 1 gnd
rlabel metal1 -26 -414 -15 -410 5 vdd
rlabel metal1 -29 -509 -23 -504 1 gnd
rlabel metal1 122 -424 126 -419 1 c4
rlabel metal1 -168 305 -164 309 5 vdd
rlabel metal1 -119 198 -113 202 1 gnd
rlabel metal1 -76 244 -70 248 1 gnd
rlabel metal1 -176 244 -170 247 1 gnd
rlabel metal1 -76 305 -71 309 5 vdd
rlabel metal1 -139 305 -134 309 5 vdd
rlabel metal1 71 139 75 143 5 vdd
rlabel metal1 120 32 126 36 1 gnd
rlabel metal1 163 78 169 82 1 gnd
rlabel metal1 63 78 69 81 1 gnd
rlabel metal1 163 139 168 143 5 vdd
rlabel metal1 100 139 105 143 5 vdd
rlabel metal1 131 -22 135 -18 5 vdd
rlabel metal1 180 -129 186 -125 1 gnd
rlabel metal1 223 -83 229 -79 1 gnd
rlabel metal1 123 -83 129 -80 1 gnd
rlabel metal1 223 -22 228 -18 5 vdd
rlabel metal1 160 -22 165 -18 5 vdd
rlabel metal2 -54 245 -50 251 1 sum1
rlabel metal2 185 79 189 85 1 sum2
rlabel metal2 245 -82 249 -76 7 sum3
rlabel metal1 -709 653 -705 657 3 gnd
rlabel metal1 -709 601 -705 605 3 gnd
rlabel metal1 -604 653 -600 657 3 gnd
rlabel metal1 -604 601 -600 605 3 gnd
rlabel metal1 -515 647 -512 651 7 vdd
rlabel metal1 -515 594 -512 598 7 vdd
rlabel metal1 -620 680 -617 684 3 vdd
rlabel metal1 -620 648 -617 652 3 vdd
rlabel metal1 -620 593 -617 597 3 vdd
rlabel metal1 -684 681 -681 684 3 gnd
rlabel metal1 -709 445 -705 449 3 gnd
rlabel metal1 -709 393 -705 397 3 gnd
rlabel metal1 -604 445 -600 449 3 gnd
rlabel metal1 -604 393 -600 397 3 gnd
rlabel metal1 -515 439 -512 443 7 vdd
rlabel metal1 -515 386 -512 390 7 vdd
rlabel metal1 -620 472 -617 476 3 vdd
rlabel metal1 -620 440 -617 444 3 vdd
rlabel metal1 -620 385 -617 389 3 vdd
rlabel metal1 -684 473 -681 476 3 gnd
rlabel metal1 -530 738 -527 742 3 vdd
rlabel metal1 -594 739 -591 742 3 gnd
rlabel metal1 -448 677 -444 681 3 gnd
rlabel metal1 -448 625 -444 629 3 gnd
rlabel metal1 -343 677 -339 681 3 gnd
rlabel metal1 -343 625 -339 629 3 gnd
rlabel metal1 -254 671 -251 675 7 vdd
rlabel metal1 -254 618 -251 622 7 vdd
rlabel metal1 -359 704 -356 708 3 vdd
rlabel metal1 -359 672 -356 676 3 vdd
rlabel metal1 -359 617 -356 621 3 vdd
rlabel metal1 -423 705 -420 708 3 gnd
rlabel metal1 -448 469 -444 473 3 gnd
rlabel metal1 -448 417 -444 421 3 gnd
rlabel metal1 -343 469 -339 473 3 gnd
rlabel metal1 -343 417 -339 421 3 gnd
rlabel metal1 -254 463 -251 467 7 vdd
rlabel metal1 -254 410 -251 414 7 vdd
rlabel metal1 -359 496 -356 500 3 vdd
rlabel metal1 -359 464 -356 468 3 vdd
rlabel metal1 -359 409 -356 413 3 vdd
rlabel metal1 -423 497 -420 500 3 gnd
rlabel metal1 -269 762 -266 766 3 vdd
rlabel metal1 -333 763 -330 766 3 gnd
rlabel metal1 -737 111 -733 115 1 gnd
rlabel metal1 -685 111 -681 115 1 gnd
rlabel metal1 -737 216 -733 220 1 gnd
rlabel metal1 -685 216 -681 220 1 gnd
rlabel metal1 -731 305 -727 308 5 vdd
rlabel metal1 -678 305 -674 308 5 vdd
rlabel metal1 -764 200 -760 203 1 vdd
rlabel metal1 -732 200 -728 203 1 vdd
rlabel metal1 -677 200 -673 203 1 vdd
rlabel metal1 -764 136 -761 139 1 gnd
rlabel metal1 -529 111 -525 115 1 gnd
rlabel metal1 -477 111 -473 115 1 gnd
rlabel metal1 -529 216 -525 220 1 gnd
rlabel metal1 -477 216 -473 220 1 gnd
rlabel metal1 -523 305 -519 308 5 vdd
rlabel metal1 -470 305 -466 308 5 vdd
rlabel metal1 -556 200 -552 203 1 vdd
rlabel metal1 -524 200 -520 203 1 vdd
rlabel metal1 -469 200 -465 203 1 vdd
rlabel metal1 -556 136 -553 139 1 gnd
rlabel metal1 -822 290 -818 293 1 vdd
rlabel metal1 -822 226 -819 229 1 gnd
rlabel metal1 -954 662 -950 666 3 gnd
rlabel metal1 -954 610 -950 614 3 gnd
rlabel metal1 -849 662 -845 666 3 gnd
rlabel metal1 -849 610 -845 614 3 gnd
rlabel metal1 -760 656 -757 660 7 vdd
rlabel metal1 -760 603 -757 607 7 vdd
rlabel metal1 -865 689 -862 693 3 vdd
rlabel metal1 -865 657 -862 661 3 vdd
rlabel metal1 -865 602 -862 606 3 vdd
rlabel metal1 -929 690 -926 693 3 gnd
rlabel metal1 -954 454 -950 458 3 gnd
rlabel metal1 -954 402 -950 406 3 gnd
rlabel metal1 -849 454 -845 458 3 gnd
rlabel metal1 -849 402 -845 406 3 gnd
rlabel metal1 -760 448 -757 452 7 vdd
rlabel metal1 -760 395 -757 399 7 vdd
rlabel metal1 -865 481 -862 485 3 vdd
rlabel metal1 -865 449 -862 453 3 vdd
rlabel metal1 -865 394 -862 398 3 vdd
rlabel metal1 -929 482 -926 485 3 gnd
rlabel metal1 -775 747 -772 751 3 vdd
rlabel metal1 -839 748 -836 751 3 gnd
rlabel metal1 -750 -103 -746 -99 1 gnd
rlabel metal1 -698 -103 -694 -99 1 gnd
rlabel metal1 -750 2 -746 6 1 gnd
rlabel metal1 -698 2 -694 6 1 gnd
rlabel metal1 -744 91 -740 94 5 vdd
rlabel metal1 -691 91 -687 94 5 vdd
rlabel metal1 -777 -14 -773 -11 1 vdd
rlabel metal1 -745 -14 -741 -11 1 vdd
rlabel metal1 -690 -14 -686 -11 1 vdd
rlabel metal1 -777 -78 -774 -75 1 gnd
rlabel metal1 -542 -103 -538 -99 1 gnd
rlabel metal1 -490 -103 -486 -99 1 gnd
rlabel metal1 -542 2 -538 6 1 gnd
rlabel metal1 -490 2 -486 6 1 gnd
rlabel metal1 -536 91 -532 94 5 vdd
rlabel metal1 -483 91 -479 94 5 vdd
rlabel metal1 -569 -14 -565 -11 1 vdd
rlabel metal1 -537 -14 -533 -11 1 vdd
rlabel metal1 -482 -14 -478 -11 1 vdd
rlabel metal1 -569 -78 -566 -75 1 gnd
rlabel metal1 -835 76 -831 79 1 vdd
rlabel metal1 -835 12 -832 15 1 gnd
rlabel metal1 -957 301 -954 304 3 gnd
rlabel metal1 -893 300 -890 304 3 vdd
rlabel metal1 -1047 35 -1044 38 3 gnd
rlabel metal1 -983 -53 -980 -49 3 vdd
rlabel metal1 -983 2 -980 6 3 vdd
rlabel metal1 -983 34 -980 38 3 vdd
rlabel metal1 -878 -52 -875 -48 7 vdd
rlabel metal1 -878 1 -875 5 7 vdd
rlabel metal1 -967 -45 -963 -41 3 gnd
rlabel metal1 -967 7 -963 11 3 gnd
rlabel metal1 -1072 -45 -1068 -41 3 gnd
rlabel metal1 -1072 7 -1068 11 3 gnd
rlabel metal1 -1047 243 -1044 246 3 gnd
rlabel metal1 -983 155 -980 159 3 vdd
rlabel metal1 -983 210 -980 214 3 vdd
rlabel metal1 -983 242 -980 246 3 vdd
rlabel metal1 -878 156 -875 160 7 vdd
rlabel metal1 -878 209 -875 213 7 vdd
rlabel metal1 -967 163 -963 167 3 gnd
rlabel metal1 -967 215 -963 219 3 gnd
rlabel metal1 -1072 163 -1068 167 3 gnd
rlabel metal1 -1072 215 -1068 219 3 gnd
rlabel metal1 -837 -219 -834 -216 1 gnd
rlabel metal1 -837 -155 -833 -152 1 vdd
rlabel metal1 -571 -309 -568 -306 1 gnd
rlabel metal1 -484 -245 -480 -242 1 vdd
rlabel metal1 -539 -245 -535 -242 1 vdd
rlabel metal1 -571 -245 -567 -242 1 vdd
rlabel metal1 -485 -140 -481 -137 5 vdd
rlabel metal1 -538 -140 -534 -137 5 vdd
rlabel metal1 -492 -229 -488 -225 1 gnd
rlabel metal1 -544 -229 -540 -225 1 gnd
rlabel metal1 -492 -334 -488 -330 1 gnd
rlabel metal1 -544 -334 -540 -330 1 gnd
rlabel metal1 -779 -309 -776 -306 1 gnd
rlabel metal1 -692 -245 -688 -242 1 vdd
rlabel metal1 -747 -245 -743 -242 1 vdd
rlabel metal1 -779 -245 -775 -242 1 vdd
rlabel metal1 -693 -140 -689 -137 5 vdd
rlabel metal1 -746 -140 -742 -137 5 vdd
rlabel metal1 -700 -229 -696 -225 1 gnd
rlabel metal1 -752 -229 -748 -225 1 gnd
rlabel metal1 -700 -334 -696 -330 1 gnd
rlabel metal1 -752 -334 -748 -330 1 gnd
rlabel metal1 -846 -434 -843 -431 1 gnd
rlabel metal1 -846 -370 -842 -367 1 vdd
rlabel metal1 -580 -524 -577 -521 1 gnd
rlabel metal1 -493 -460 -489 -457 1 vdd
rlabel metal1 -548 -460 -544 -457 1 vdd
rlabel metal1 -580 -460 -576 -457 1 vdd
rlabel metal1 -494 -355 -490 -352 5 vdd
rlabel metal1 -547 -355 -543 -352 5 vdd
rlabel metal1 -501 -444 -497 -440 1 gnd
rlabel metal1 -553 -444 -549 -440 1 gnd
rlabel metal1 -501 -549 -497 -545 1 gnd
rlabel metal1 -553 -549 -549 -545 1 gnd
rlabel metal1 -788 -524 -785 -521 1 gnd
rlabel metal1 -701 -460 -697 -457 1 vdd
rlabel metal1 -756 -460 -752 -457 1 vdd
rlabel metal1 -788 -460 -784 -457 1 vdd
rlabel metal1 -702 -355 -698 -352 5 vdd
rlabel metal1 -755 -355 -751 -352 5 vdd
rlabel metal1 -709 -444 -705 -440 1 gnd
rlabel metal1 -761 -444 -757 -440 1 gnd
rlabel metal1 -709 -549 -705 -545 1 gnd
rlabel metal1 -761 -549 -757 -545 1 gnd
rlabel metal1 -200 486 -197 489 1 gnd
rlabel metal1 -200 550 -196 553 1 vdd
rlabel metal1 66 396 69 399 1 gnd
rlabel metal1 153 460 157 463 1 vdd
rlabel metal1 98 460 102 463 1 vdd
rlabel metal1 66 460 70 463 1 vdd
rlabel metal1 152 565 156 568 5 vdd
rlabel metal1 99 565 103 568 5 vdd
rlabel metal1 145 476 149 480 1 gnd
rlabel metal1 93 476 97 480 1 gnd
rlabel metal1 145 371 149 375 1 gnd
rlabel metal1 93 371 97 375 1 gnd
rlabel metal1 -142 396 -139 399 1 gnd
rlabel metal1 -55 460 -51 463 1 vdd
rlabel metal1 -110 460 -106 463 1 vdd
rlabel metal1 -142 460 -138 463 1 vdd
rlabel metal1 -56 565 -52 568 5 vdd
rlabel metal1 -109 565 -105 568 5 vdd
rlabel metal1 -63 476 -59 480 1 gnd
rlabel metal1 -115 476 -111 480 1 gnd
rlabel metal1 -63 371 -59 375 1 gnd
rlabel metal1 -115 371 -111 375 1 gnd
rlabel metal1 74 281 77 284 1 gnd
rlabel metal1 74 345 78 348 1 vdd
rlabel metal1 340 191 343 194 1 gnd
rlabel metal1 427 255 431 258 1 vdd
rlabel metal1 372 255 376 258 1 vdd
rlabel metal1 340 255 344 258 1 vdd
rlabel metal1 426 360 430 363 5 vdd
rlabel metal1 373 360 377 363 5 vdd
rlabel metal1 419 271 423 275 1 gnd
rlabel metal1 367 271 371 275 1 gnd
rlabel metal1 419 166 423 170 1 gnd
rlabel metal1 367 166 371 170 1 gnd
rlabel metal1 132 191 135 194 1 gnd
rlabel metal1 219 255 223 258 1 vdd
rlabel metal1 164 255 168 258 1 vdd
rlabel metal1 132 255 136 258 1 vdd
rlabel metal1 218 360 222 363 5 vdd
rlabel metal1 165 360 169 363 5 vdd
rlabel metal1 211 271 215 275 1 gnd
rlabel metal1 159 271 163 275 1 gnd
rlabel metal1 211 166 215 170 1 gnd
rlabel metal1 159 166 163 170 1 gnd
rlabel metal1 380 -61 384 -57 1 gnd
rlabel metal1 432 -61 436 -57 1 gnd
rlabel metal1 380 44 384 48 1 gnd
rlabel metal1 432 44 436 48 1 gnd
rlabel metal1 386 133 390 136 5 vdd
rlabel metal1 439 133 443 136 5 vdd
rlabel metal1 353 28 357 31 1 vdd
rlabel metal1 385 28 389 31 1 vdd
rlabel metal1 440 28 444 31 1 vdd
rlabel metal1 353 -36 356 -33 1 gnd
rlabel metal1 588 -61 592 -57 1 gnd
rlabel metal1 640 -61 644 -57 1 gnd
rlabel metal1 588 44 592 48 1 gnd
rlabel metal1 640 44 644 48 1 gnd
rlabel metal1 594 133 598 136 5 vdd
rlabel metal1 647 133 651 136 5 vdd
rlabel metal1 561 28 565 31 1 vdd
rlabel metal1 593 28 597 31 1 vdd
rlabel metal1 648 28 652 31 1 vdd
rlabel metal1 561 -36 564 -33 1 gnd
rlabel metal1 295 118 299 121 1 vdd
rlabel metal1 295 54 298 57 1 gnd
rlabel metal1 374 -275 378 -271 1 gnd
rlabel metal1 426 -275 430 -271 1 gnd
rlabel metal1 374 -170 378 -166 1 gnd
rlabel metal1 426 -170 430 -166 1 gnd
rlabel metal1 380 -81 384 -78 5 vdd
rlabel metal1 433 -81 437 -78 5 vdd
rlabel metal1 347 -186 351 -183 1 vdd
rlabel metal1 379 -186 383 -183 1 vdd
rlabel metal1 434 -186 438 -183 1 vdd
rlabel metal1 347 -250 350 -247 1 gnd
rlabel metal1 582 -275 586 -271 1 gnd
rlabel metal1 634 -275 638 -271 1 gnd
rlabel metal1 582 -170 586 -166 1 gnd
rlabel metal1 634 -170 638 -166 1 gnd
rlabel metal1 588 -81 592 -78 5 vdd
rlabel metal1 641 -81 645 -78 5 vdd
rlabel metal1 555 -186 559 -183 1 vdd
rlabel metal1 587 -186 591 -183 1 vdd
rlabel metal1 642 -186 646 -183 1 vdd
rlabel metal1 555 -250 558 -247 1 gnd
rlabel metal1 289 -96 293 -93 1 vdd
rlabel metal1 289 -160 292 -157 1 gnd
rlabel metal1 287 -499 291 -495 1 gnd
rlabel metal1 339 -499 343 -495 1 gnd
rlabel metal1 287 -394 291 -390 1 gnd
rlabel metal1 339 -394 343 -390 1 gnd
rlabel metal1 293 -305 297 -302 5 vdd
rlabel metal1 346 -305 350 -302 5 vdd
rlabel metal1 260 -410 264 -407 1 vdd
rlabel metal1 292 -410 296 -407 1 vdd
rlabel metal1 347 -410 351 -407 1 vdd
rlabel metal1 260 -474 263 -471 1 gnd
rlabel metal1 495 -499 499 -495 1 gnd
rlabel metal1 547 -499 551 -495 1 gnd
rlabel metal1 495 -394 499 -390 1 gnd
rlabel metal1 547 -394 551 -390 1 gnd
rlabel metal1 501 -305 505 -302 5 vdd
rlabel metal1 554 -305 558 -302 5 vdd
rlabel metal1 468 -410 472 -407 1 vdd
rlabel metal1 500 -410 504 -407 1 vdd
rlabel metal1 555 -410 559 -407 1 vdd
rlabel metal1 468 -474 471 -471 1 gnd
rlabel metal1 202 -320 206 -317 1 vdd
rlabel metal1 202 -384 205 -381 1 gnd
rlabel metal1 -812 -403 -809 -398 1 bin_3
rlabel metal1 -803 -188 -800 -183 1 ain_3
rlabel metal1 -926 265 -921 270 1 bin_2
rlabel metal1 -798 43 -793 48 1 ain_2
rlabel metal1 -789 257 -784 262 1 bin_1
rlabel metal1 -808 711 -803 716 1 ain_1
rlabel metal1 -563 703 -558 708 1 bin_0
rlabel metal1 -302 727 -297 732 1 ain_0
rlabel metal1 199 514 205 518 1 sumo_0
rlabel metal1 474 309 478 313 1 sumo_1
rlabel metal1 701 82 706 86 7 sumo_2
rlabel metal1 689 -132 693 -128 1 sumo_3
rlabel metal1 601 -356 605 -352 1 c_out
rlabel metal1 -898 777 -892 781 1 clk
<< end >>
