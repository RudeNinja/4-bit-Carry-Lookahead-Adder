* SPICE3 file created from carry.ext - technology: scmos

.option scale=0.09u
.include TSMC_180nm.txt
.param SUPPLY=1.8

.global gnd vdd
Vdd vdd gnd 'SUPPLY'


vin_a1 Pi gnd  pulse 0 1.8 0ns 100ps 100ps 4.9ns 10ns
vin_a2 Cin gnd pulse 0 1.8 0ns 100ps 100ps 9.9ns 20ns
vin_a3 Gi gnd pulse 0 1.8 0ns 100ps 100ps 19.9ns 40ns

M1000 a_n37_n13# Pi gnd Gnd CMOSN w=8 l=2
+  ad=88 pd=38 as=264 ps=146
M1001 a_66_35# Gi vdd Vdd CMOSP w=11 l=2
+  ad=176 pd=54 as=462 ps=194
M1002 a_n37_36# Cin a_n37_n13# Gnd CMOSN w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1003 a_66_n26# a_n2_n12# a_66_35# Vdd CMOSP w=11 l=2
+  ad=99 pd=40 as=0 ps=0
M1004 a_n2_n12# a_n37_36# gnd Gnd CMOSN w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1005 C_out a_66_n26# gnd Gnd CMOSN w=8 l=2
+  ad=56 pd=30 as=0 ps=0
M1006 vdd Cin a_n37_36# Vdd CMOSP w=11 l=2
+  ad=0 pd=0 as=121 ps=44
M1007 a_n37_36# Pi vdd Vdd CMOSP w=11 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 gnd a_n2_n12# a_66_n26# Gnd CMOSN w=8 l=2
+  ad=0 pd=0 as=128 ps=48
M1009 C_out a_66_n26# vdd Vdd CMOSP w=11 l=2
+  ad=99 pd=40 as=0 ps=0
M1010 a_66_n26# Gi gnd Gnd CMOSN w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 a_n2_n12# a_n37_36# vdd Vdd CMOSP w=11 l=2
+  ad=66 pd=34 as=0 ps=0
C0 a_66_n26# gnd 0.07fF
C1 a_n37_36# vdd 0.09fF
C2 a_n2_n12# a_66_n26# 0.12fF
C3 a_n37_36# gnd 0.03fF
C4 a_n37_36# a_n2_n12# 0.04fF
C5 a_66_n26# Vdd 0.12fF
C6 vdd Vdd 0.11fF
C7 a_n2_n12# Vdd 0.03fF
C8 a_n2_n12# gnd 0.07fF
C9 a_66_n26# C_out 0.04fF
C10 vdd Vdd 0.08fF
C11 a_n2_n12# Vdd 0.08fF
C12 Pi Cin 0.01fF
C13 Vdd Pi 0.06fF
C14 C_out gnd 0.05fF
C15 a_n2_n12# Gi 0.06fF
C16 Gi Vdd 0.08fF
C17 a_n37_36# Cin 0.13fF
C18 C_out Vdd 0.03fF
C19 a_n37_36# Vdd 0.09fF
C20 Vdd Cin 0.06fF
C21 gnd Gnd 0.44fF
C22 C_out Gnd 0.17fF
C23 vdd Gnd 0.33fF
C24 a_66_n26# Gnd 0.59fF
C25 Gi Gnd 0.37fF
C26 a_n2_n12# Gnd 0.71fF
C27 a_n37_36# Gnd 0.17fF
C28 Cin Gnd 0.29fF
C29 Pi Gnd 0.29fF
C30 Vdd Gnd 2.25fF
C31 Vdd Gnd 1.43fF

.control
set hcopypscolor = 1 *White background for saving plots
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7))
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7))

tran 0.1n 200n
set curplottitle= ShubhamPriyadarshan-2020102027_Q5

plot v(Pi)+2 v(Cin)+4 v(Gi)+6 v(C_out)

hardcopy Carry.ps v(Pi)+2 v(Cin)+4 v(Gi)+6 v(C_out)


.endc
.end
